
module prime_DW_mult_uns_0 ( a, b, product );
  input [10:0] a;
  input [10:0] b;
  output [21:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n40, n42, n43, n45, n46, n47, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, \a[0] , n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120;
  assign product[0] = \a[0] ;
  assign \a[0]  = a[0];

  FA1A U3 ( .A(n15), .B(n20), .CI(n3), .CO(n2), .S(product[9]) );
  FA1A U4 ( .A(n21), .B(n26), .CI(n4), .CO(n3), .S(product[8]) );
  FA1A U7 ( .A(n35), .B(n36), .CI(n7), .CO(n6), .S(product[5]) );
  FA1A U8 ( .A(n37), .B(n59), .CI(n8), .CO(n7), .S(product[4]) );
  HA1 U9 ( .A(n9), .B(n61), .CO(n8), .S(product[3]) );
  HA1 U10 ( .A(n62), .B(a[1]), .CO(n9), .S(product[2]) );
  FA1A U15 ( .A(n22), .B(n19), .CI(n17), .CO(n14), .S(n15) );
  FA1A U16 ( .A(n45), .B(n49), .CI(n24), .CO(n16), .S(n17) );
  HA1 U17 ( .A(n40), .B(n42), .CO(n18), .S(n19) );
  FA1A U18 ( .A(n25), .B(n50), .CI(n23), .CO(n20), .S(n21) );
  FA1A U19 ( .A(n43), .B(n53), .CI(n28), .CO(n22), .S(n23) );
  FA1A U21 ( .A(n32), .B(n51), .CI(n29), .CO(n26), .S(n27) );
  HA1 U22 ( .A(n47), .B(n54), .CO(n28), .S(n29) );
  FA1A U23 ( .A(n52), .B(n55), .CI(n34), .CO(n30), .S(n31) );
  HA1 U25 ( .A(n56), .B(n58), .CO(n34), .S(n35) );
  HA1 U26 ( .A(n60), .B(a[2]), .CO(n36), .S(n37) );
  IV U68 ( .A(b[1]), .Z(n100) );
  FA1AP U69 ( .A(n27), .B(n30), .CI(n5), .CO(n4), .S(product[7]) );
  IVP U70 ( .A(b[5]), .Z(n105) );
  FA1A U71 ( .A(n31), .B(n33), .CI(n6), .CO(n5), .S(product[6]) );
  HA1 U72 ( .A(n46), .B(a[4]), .CO(n24), .S(n25) );
  IVDA U73 ( .A(b[6]), .Y(n106) );
  IVDA U74 ( .A(b[7]), .Y(n107) );
  HA1 U75 ( .A(n57), .B(a[3]), .CO(n32), .S(n33) );
  IV U76 ( .A(b[4]), .Z(n104) );
  IV U77 ( .A(b[3]), .Z(n103) );
  IV U78 ( .A(b[2]), .Z(n102) );
  IV U79 ( .A(b[0]), .Z(n101) );
  EO U80 ( .A(n108), .B(n109), .Z(product[10]) );
  EN U81 ( .A(n2), .B(n14), .Z(n109) );
  EO U82 ( .A(n110), .B(n111), .Z(n108) );
  EO U83 ( .A(n112), .B(n113), .Z(n111) );
  EO U84 ( .A(n114), .B(n115), .Z(n113) );
  ND2 U85 ( .A(b[0]), .B(b[9]), .Z(n115) );
  ND2 U86 ( .A(b[4]), .B(b[5]), .Z(n114) );
  EO U87 ( .A(n116), .B(n117), .Z(n112) );
  ND2 U88 ( .A(b[2]), .B(b[7]), .Z(n117) );
  ND2 U89 ( .A(b[3]), .B(b[6]), .Z(n116) );
  EO U90 ( .A(n118), .B(n119), .Z(n110) );
  EN U91 ( .A(n105), .B(n18), .Z(n119) );
  EO U92 ( .A(n120), .B(n16), .Z(n118) );
  ND2 U93 ( .A(b[1]), .B(b[8]), .Z(n120) );
  NR2 U94 ( .A(n100), .B(n101), .Z(n62) );
  NR2 U95 ( .A(n102), .B(n101), .Z(n61) );
  NR2 U96 ( .A(n100), .B(n102), .Z(n60) );
  NR2 U97 ( .A(n103), .B(n101), .Z(n59) );
  NR2 U98 ( .A(n100), .B(n103), .Z(n58) );
  NR2 U99 ( .A(n103), .B(n102), .Z(n57) );
  NR2 U100 ( .A(n104), .B(n101), .Z(n56) );
  NR2 U101 ( .A(n100), .B(n104), .Z(n55) );
  NR2 U102 ( .A(n102), .B(n104), .Z(n54) );
  NR2 U103 ( .A(n103), .B(n104), .Z(n53) );
  NR2 U104 ( .A(n105), .B(n101), .Z(n52) );
  NR2 U105 ( .A(n105), .B(n100), .Z(n51) );
  NR2 U106 ( .A(n105), .B(n102), .Z(n50) );
  NR2 U107 ( .A(n105), .B(n103), .Z(n49) );
  NR2 U108 ( .A(n106), .B(n101), .Z(n47) );
  NR2 U109 ( .A(n100), .B(n106), .Z(n46) );
  NR2 U110 ( .A(n106), .B(n102), .Z(n45) );
  NR2 U111 ( .A(n107), .B(n101), .Z(n43) );
  NR2 U112 ( .A(n100), .B(n107), .Z(n42) );
  AN2 U113 ( .A(b[8]), .B(b[0]), .Z(n40) );
endmodule


module prime_DW01_add_25 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , \A[1] , n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];

  ND4 U36 ( .A(n81), .B(n72), .C(n88), .D(n89), .Z(n83) );
  ND2 U37 ( .A(A[5]), .B(B[5]), .Z(n85) );
  ND2 U38 ( .A(A[5]), .B(B[5]), .Z(n72) );
  ND2 U39 ( .A(n88), .B(n89), .Z(n80) );
  IVDA U40 ( .A(B[4]), .Y(n69), .Z(n70) );
  B2I U41 ( .A(B[3]), .Z2(n71) );
  EOP U42 ( .A(n74), .B(n73), .Z(n79) );
  NR2P U43 ( .A(n70), .B(A[4]), .Z(n74) );
  NR2P U44 ( .A(A[5]), .B(B[5]), .Z(n86) );
  AO1P U45 ( .A(n74), .B(n85), .C(n86), .D(n87), .Z(n84) );
  EOP U46 ( .A(A[5]), .B(B[5]), .Z(n73) );
  EO U47 ( .A(n81), .B(n73), .Z(n78) );
  EO U48 ( .A(n77), .B(B[2]), .Z(SUM[2]) );
  MUX21L U49 ( .A(n78), .B(n79), .S(n80), .Z(SUM[5]) );
  EO3 U50 ( .A(A[3]), .B(n71), .C(n82), .Z(SUM[3]) );
  EO3 U51 ( .A(A[4]), .B(n75), .C(n80), .Z(SUM[4]) );
  ND2 U52 ( .A(A[3]), .B(n71), .Z(n89) );
  IVA U53 ( .A(n69), .Z(n75) );
  IV U54 ( .A(B[2]), .Z(n76) );
  IVA U55 ( .A(A[2]), .Z(n77) );
  AN2P U56 ( .A(n83), .B(n84), .Z(CO) );
  ND8 U57 ( .A(B[6]), .B(B[7]), .C(B[13]), .D(B[9]), .E(B[8]), .F(B[11]), .G(
        B[10]), .H(B[12]), .Z(n87) );
  AO7P U58 ( .A(A[3]), .B(n71), .C(n82), .Z(n88) );
  ND2P U59 ( .A(n76), .B(n77), .Z(n82) );
  ND2P U60 ( .A(n75), .B(A[4]), .Z(n81) );
endmodule


module prime_DW01_add_74 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n33, n34, n35, n36,
         n37, n38, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n64, n65, n66, n67, n68, n69,
         n70, \A[0] , n118, n119, n120, n121, n122, n123;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  NR2 U7 ( .A(n18), .B(n16), .Z(n14) );
  NR2 U9 ( .A(A[11]), .B(B[11]), .Z(n16) );
  NR2 U11 ( .A(A[10]), .B(B[10]), .Z(n18) );
  NR2 U25 ( .A(n37), .B(n30), .Z(n28) );
  NR2 U39 ( .A(n41), .B(n46), .Z(n35) );
  NR2 U51 ( .A(A[6]), .B(B[6]), .Z(n46) );
  NR2 U56 ( .A(n55), .B(n52), .Z(n50) );
  FA1A U76 ( .A(B[2]), .B(A[2]), .CI(n123), .CO(n61), .S(SUM[2]) );
  IV U84 ( .A(n69), .Z(n118) );
  AO7P U85 ( .A(n41), .B(n47), .C(n42), .Z(n36) );
  ND2P U86 ( .A(A[4]), .B(B[4]), .Z(n56) );
  AO6 U87 ( .A(n50), .B(n58), .C(n51), .Z(n49) );
  AN2 U88 ( .A(n15), .B(B[12]), .Z(n119) );
  AN2 U89 ( .A(n14), .B(B[12]), .Z(n120) );
  NR2P U90 ( .A(n25), .B(n30), .Z(n23) );
  AO7 U91 ( .A(n121), .B(n21), .C(n22), .Z(n20) );
  ENP U92 ( .A(n8), .B(n61), .Z(SUM[3]) );
  AO6 U93 ( .A(n23), .B(n36), .C(n24), .Z(n22) );
  NR2P U94 ( .A(A[7]), .B(B[7]), .Z(n41) );
  AO6 U95 ( .A(n122), .B(n35), .C(n36), .Z(n34) );
  NR2P U96 ( .A(A[9]), .B(B[9]), .Z(n25) );
  AO6P U97 ( .A(n50), .B(n58), .C(n51), .Z(n121) );
  AO7P U98 ( .A(n59), .B(n1), .C(n60), .Z(n58) );
  NR2P U99 ( .A(A[4]), .B(B[4]), .Z(n55) );
  IV U100 ( .A(n49), .Z(n122) );
  NR2P U101 ( .A(A[3]), .B(B[3]), .Z(n59) );
  AO7P U102 ( .A(n52), .B(n56), .C(n53), .Z(n51) );
  NR2P U103 ( .A(A[8]), .B(B[8]), .Z(n30) );
  EOP U104 ( .A(n34), .B(n3), .Z(SUM[8]) );
  IVP U105 ( .A(n9), .Z(CO) );
  IV U106 ( .A(n41), .Z(n66) );
  IV U107 ( .A(n47), .Z(n45) );
  AO6P U108 ( .A(n20), .B(n120), .C(n119), .Z(n9) );
  IV U109 ( .A(n58), .Z(n57) );
  ND2 U110 ( .A(n35), .B(n23), .Z(n21) );
  AO7 U111 ( .A(n25), .B(n33), .C(n26), .Z(n24) );
  IV U112 ( .A(n35), .Z(n37) );
  ND2 U113 ( .A(n65), .B(n33), .Z(n3) );
  EO U114 ( .A(n27), .B(n2), .Z(SUM[9]) );
  ND2 U115 ( .A(n64), .B(n26), .Z(n2) );
  IV U116 ( .A(n25), .Z(n64) );
  IV U117 ( .A(n36), .Z(n38) );
  ND2 U118 ( .A(A[7]), .B(B[7]), .Z(n42) );
  EN U119 ( .A(n48), .B(n5), .Z(SUM[6]) );
  ND2 U120 ( .A(n67), .B(n47), .Z(n5) );
  IV U121 ( .A(n46), .Z(n67) );
  ND2 U122 ( .A(A[6]), .B(B[6]), .Z(n47) );
  ND2 U123 ( .A(A[8]), .B(B[8]), .Z(n33) );
  ND2 U124 ( .A(A[9]), .B(B[9]), .Z(n26) );
  EN U125 ( .A(n54), .B(n6), .Z(SUM[5]) );
  ND2 U126 ( .A(n68), .B(n53), .Z(n6) );
  IV U127 ( .A(n52), .Z(n68) );
  EO U128 ( .A(n7), .B(n57), .Z(SUM[4]) );
  ND2 U129 ( .A(n69), .B(n56), .Z(n7) );
  IVP U130 ( .A(n61), .Z(n1) );
  AO7 U131 ( .A(n16), .B(n19), .C(n17), .Z(n15) );
  ND2 U132 ( .A(A[10]), .B(B[10]), .Z(n19) );
  ND2 U133 ( .A(n70), .B(n60), .Z(n8) );
  IV U134 ( .A(n59), .Z(n70) );
  EO U135 ( .A(n43), .B(n4), .Z(SUM[7]) );
  ND2 U136 ( .A(n66), .B(n42), .Z(n4) );
  OR2 U137 ( .A(B[1]), .B(A[1]), .Z(n123) );
  EN U138 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  AO7 U139 ( .A(n38), .B(n30), .C(n33), .Z(n29) );
  IV U140 ( .A(n30), .Z(n65) );
  IV U141 ( .A(n55), .Z(n69) );
  ND2 U142 ( .A(A[11]), .B(B[11]), .Z(n17) );
  IV U143 ( .A(n121), .Z(n48) );
  AO6 U144 ( .A(n28), .B(n48), .C(n29), .Z(n27) );
  AO6 U145 ( .A(n48), .B(n67), .C(n45), .Z(n43) );
  ND2 U146 ( .A(A[5]), .B(B[5]), .Z(n53) );
  AO7 U147 ( .A(n57), .B(n118), .C(n56), .Z(n54) );
  ND2 U148 ( .A(A[3]), .B(B[3]), .Z(n60) );
  NR2P U149 ( .A(A[5]), .B(B[5]), .Z(n52) );
endmodule


module prime_DW01_add_88 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n51, n52, n53,
         n54, n56, n103, n104, n105, n106;

  NR2 U4 ( .A(n24), .B(n104), .Z(n12) );
  NR2 U5 ( .A(n25), .B(n104), .Z(n13) );
  NR2 U10 ( .A(n20), .B(n19), .Z(n18) );
  NR2 U13 ( .A(n23), .B(n22), .Z(n21) );
  NR2 U19 ( .A(A[8]), .B(B[8]), .Z(n24) );
  NR2 U29 ( .A(A[7]), .B(B[7]), .Z(n31) );
  MUX21LP U38 ( .A(n38), .B(n37), .S(n45), .Z(n36) );
  NR2 U57 ( .A(A[3]), .B(B[3]), .Z(n46) );
  FA1A U59 ( .A(n49), .B(A[2]), .CI(B[2]), .CO(n48), .S(SUM[2]) );
  FA1A U60 ( .A(n106), .B(A[1]), .CI(B[1]), .CO(n49), .S(SUM[1]) );
  MUX21L U68 ( .A(n10), .B(n11), .S(n36), .Z(CO) );
  NR2P U69 ( .A(A[5]), .B(B[5]), .Z(n39) );
  MUX21LP U70 ( .A(n31), .B(n32), .S(n35), .Z(n30) );
  IVAP U71 ( .A(n103), .Z(n42) );
  EOP U72 ( .A(n36), .B(n5), .Z(SUM[6]) );
  OR2P U73 ( .A(A[4]), .B(B[4]), .Z(n103) );
  MUX21LP U74 ( .A(n31), .B(n32), .S(n34), .Z(n29) );
  NR2P U75 ( .A(A[6]), .B(B[6]), .Z(n34) );
  ENP U76 ( .A(n41), .B(n6), .Z(SUM[5]) );
  ENP U77 ( .A(n26), .B(n3), .Z(SUM[8]) );
  IV U78 ( .A(B[10]), .Z(n23) );
  IV U79 ( .A(B[12]), .Z(n19) );
  IV U80 ( .A(B[11]), .Z(n22) );
  AN2 U81 ( .A(n18), .B(B[13]), .Z(n105) );
  MUX21LP U82 ( .A(n47), .B(n46), .S(n48), .Z(n45) );
  ND2 U83 ( .A(n103), .B(n43), .Z(n7) );
  EN U84 ( .A(n33), .B(n4), .Z(SUM[7]) );
  ND2 U85 ( .A(n52), .B(n32), .Z(n4) );
  ND2 U86 ( .A(n54), .B(n40), .Z(n6) );
  IV U87 ( .A(n39), .Z(n54) );
  ND2 U88 ( .A(n56), .B(n47), .Z(n8) );
  ND2 U89 ( .A(n53), .B(n35), .Z(n5) );
  ND2 U90 ( .A(n51), .B(n25), .Z(n3) );
  IV U91 ( .A(n24), .Z(n51) );
  IV U92 ( .A(n31), .Z(n52) );
  EO U93 ( .A(n7), .B(n44), .Z(SUM[4]) );
  MUX21L U94 ( .A(n13), .B(n12), .S(n29), .Z(n10) );
  MUX21L U95 ( .A(n13), .B(n12), .S(n30), .Z(n11) );
  ND2 U96 ( .A(A[8]), .B(B[8]), .Z(n25) );
  MUX21H U97 ( .A(n29), .B(n30), .S(n36), .Z(n26) );
  ND2 U98 ( .A(n21), .B(B[9]), .Z(n20) );
  MUX21L U99 ( .A(n39), .B(n40), .S(n43), .Z(n38) );
  MUX21L U100 ( .A(n39), .B(n40), .S(n42), .Z(n37) );
  IVP U101 ( .A(n45), .Z(n44) );
  ND2 U102 ( .A(n105), .B(B[14]), .Z(n104) );
  EN U103 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  EN U104 ( .A(n8), .B(n48), .Z(SUM[3]) );
  OR2 U105 ( .A(B[0]), .B(A[0]), .Z(n106) );
  ND2 U106 ( .A(A[3]), .B(B[3]), .Z(n47) );
  ND2 U107 ( .A(A[6]), .B(B[6]), .Z(n35) );
  IV U108 ( .A(n46), .Z(n56) );
  MUX21L U109 ( .A(n42), .B(n43), .S(n44), .Z(n41) );
  MUX21L U110 ( .A(n34), .B(n35), .S(n36), .Z(n33) );
  IV U111 ( .A(n34), .Z(n53) );
  ND2 U112 ( .A(A[4]), .B(B[4]), .Z(n43) );
  ND2 U113 ( .A(A[5]), .B(B[5]), .Z(n40) );
  ND2 U114 ( .A(A[7]), .B(B[7]), .Z(n32) );
endmodule


module prime_DW01_add_89 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n18, n23, n24, n25, n26,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n51, n52, n56, n103, n104, n105,
         n106, n107, n108;

  NR2 U4 ( .A(n24), .B(n103), .Z(n12) );
  NR2 U5 ( .A(n25), .B(n103), .Z(n13) );
  NR2 U10 ( .A(n23), .B(n106), .Z(n18) );
  NR2 U19 ( .A(A[8]), .B(B[8]), .Z(n24) );
  NR2 U29 ( .A(A[7]), .B(B[7]), .Z(n31) );
  MUX21LP U38 ( .A(n38), .B(n37), .S(n45), .Z(n36) );
  MUX21LP U40 ( .A(n39), .B(n40), .S(n43), .Z(n38) );
  NR2 U57 ( .A(A[3]), .B(B[3]), .Z(n46) );
  FA1A U59 ( .A(n49), .B(A[2]), .CI(B[2]), .CO(n48), .S(SUM[2]) );
  FA1A U60 ( .A(n107), .B(A[1]), .CI(B[1]), .CO(n49), .S(SUM[1]) );
  ND2 U68 ( .A(n18), .B(B[13]), .Z(n103) );
  MUX21L U69 ( .A(n39), .B(n40), .S(n42), .Z(n37) );
  OR2P U70 ( .A(A[5]), .B(B[5]), .Z(n104) );
  B4I U71 ( .A(n104), .Z(n39) );
  IVAP U72 ( .A(n105), .Z(n42) );
  EOP U73 ( .A(n36), .B(n5), .Z(SUM[6]) );
  MUX21L U74 ( .A(n10), .B(n11), .S(n36), .Z(CO) );
  OR2P U75 ( .A(A[4]), .B(B[4]), .Z(n105) );
  IVAP U76 ( .A(n108), .Z(n34) );
  ENP U77 ( .A(n41), .B(n6), .Z(SUM[5]) );
  ENP U78 ( .A(n26), .B(n3), .Z(SUM[8]) );
  IV U79 ( .A(n45), .Z(n44) );
  MUX21L U80 ( .A(n13), .B(n12), .S(n30), .Z(n11) );
  MUX21L U81 ( .A(n13), .B(n12), .S(n29), .Z(n10) );
  MUX21L U82 ( .A(n31), .B(n32), .S(n35), .Z(n30) );
  MUX21L U83 ( .A(n31), .B(n32), .S(n34), .Z(n29) );
  ND2 U84 ( .A(n104), .B(n40), .Z(n6) );
  ND2 U85 ( .A(n51), .B(n25), .Z(n3) );
  EN U86 ( .A(n33), .B(n4), .Z(SUM[7]) );
  IV U87 ( .A(n24), .Z(n51) );
  ND2 U88 ( .A(n52), .B(n32), .Z(n4) );
  IV U89 ( .A(n31), .Z(n52) );
  EO U90 ( .A(n7), .B(n44), .Z(SUM[4]) );
  ND2 U91 ( .A(n105), .B(n43), .Z(n7) );
  ND2 U92 ( .A(A[8]), .B(B[8]), .Z(n25) );
  ND2 U93 ( .A(n108), .B(n35), .Z(n5) );
  MUX21H U94 ( .A(n29), .B(n30), .S(n36), .Z(n26) );
  MUX21L U95 ( .A(n34), .B(n35), .S(n36), .Z(n33) );
  ND2 U96 ( .A(B[11]), .B(B[12]), .Z(n106) );
  ND2 U97 ( .A(B[9]), .B(B[10]), .Z(n23) );
  MUX21LP U98 ( .A(n47), .B(n46), .S(n48), .Z(n45) );
  EN U99 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  EN U100 ( .A(n8), .B(n48), .Z(SUM[3]) );
  ND2 U101 ( .A(n56), .B(n47), .Z(n8) );
  OR2 U102 ( .A(B[0]), .B(A[0]), .Z(n107) );
  ND2 U103 ( .A(A[3]), .B(B[3]), .Z(n47) );
  ND2 U104 ( .A(A[6]), .B(B[6]), .Z(n35) );
  IV U105 ( .A(n46), .Z(n56) );
  MUX21L U106 ( .A(n42), .B(n43), .S(n44), .Z(n41) );
  OR2P U107 ( .A(A[6]), .B(B[6]), .Z(n108) );
  ND2 U108 ( .A(A[4]), .B(B[4]), .Z(n43) );
  ND2 U109 ( .A(A[5]), .B(B[5]), .Z(n40) );
  ND2 U110 ( .A(A[7]), .B(B[7]), .Z(n32) );
endmodule


module prime_DW01_add_87 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n19, n20, n21, n22, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n53, n54, n55,
         n56, n57, n58, n105, n106, n107, n108, n109;

  NR2 U4 ( .A(n25), .B(n107), .Z(n11) );
  NR2 U5 ( .A(n26), .B(n107), .Z(n12) );
  NR2 U12 ( .A(n21), .B(n20), .Z(n19) );
  NR2 U21 ( .A(A[8]), .B(B[8]), .Z(n25) );
  MUX21LP U28 ( .A(n32), .B(n33), .S(n36), .Z(n31) );
  NR2 U31 ( .A(A[7]), .B(B[7]), .Z(n32) );
  MUX21LP U40 ( .A(n39), .B(n38), .S(n46), .Z(n37) );
  FA1A U61 ( .A(n50), .B(A[2]), .CI(B[2]), .CO(n49), .S(SUM[2]) );
  FA1A U62 ( .A(B[1]), .B(A[1]), .CI(n109), .CO(n50), .S(SUM[1]) );
  MUX21LP U70 ( .A(n39), .B(n38), .S(n46), .Z(n105) );
  NR2 U71 ( .A(A[3]), .B(B[3]), .Z(n47) );
  EOP U72 ( .A(n105), .B(n4), .Z(SUM[6]) );
  MUX21L U73 ( .A(n40), .B(n41), .S(n43), .Z(n38) );
  NR2P U74 ( .A(A[5]), .B(B[5]), .Z(n40) );
  MUX21L U75 ( .A(n9), .B(n10), .S(n37), .Z(CO) );
  NR2P U76 ( .A(A[6]), .B(B[6]), .Z(n35) );
  NR2P U77 ( .A(A[4]), .B(B[4]), .Z(n43) );
  IV U78 ( .A(n31), .Z(n29) );
  MUX21LP U79 ( .A(n32), .B(n33), .S(n35), .Z(n30) );
  AN2P U80 ( .A(n19), .B(B[13]), .Z(n106) );
  MUX21LP U81 ( .A(n48), .B(n47), .S(n49), .Z(n46) );
  OR2P U82 ( .A(B[0]), .B(A[0]), .Z(n109) );
  IVP U83 ( .A(n30), .Z(n28) );
  MUX21L U84 ( .A(n12), .B(n11), .S(n30), .Z(n9) );
  MUX21L U85 ( .A(n12), .B(n11), .S(n31), .Z(n10) );
  ND2 U86 ( .A(A[8]), .B(B[8]), .Z(n26) );
  EN U87 ( .A(n27), .B(n2), .Z(SUM[8]) );
  ND2 U88 ( .A(n53), .B(n26), .Z(n2) );
  MUX21L U89 ( .A(n28), .B(n29), .S(n105), .Z(n27) );
  IV U90 ( .A(n25), .Z(n53) );
  EN U91 ( .A(n42), .B(n5), .Z(SUM[5]) );
  ND2 U92 ( .A(n56), .B(n41), .Z(n5) );
  IV U93 ( .A(n40), .Z(n56) );
  EN U94 ( .A(n34), .B(n3), .Z(SUM[7]) );
  ND2 U95 ( .A(n54), .B(n33), .Z(n3) );
  IV U96 ( .A(n32), .Z(n54) );
  EO U97 ( .A(n6), .B(n45), .Z(SUM[4]) );
  ND2 U98 ( .A(n57), .B(n44), .Z(n6) );
  ND2 U99 ( .A(n55), .B(n36), .Z(n4) );
  IVDA U100 ( .A(B[11]), .Y(n21) );
  IV U101 ( .A(B[12]), .Z(n20) );
  AN2P U102 ( .A(B[10]), .B(B[9]), .Z(n22) );
  MUX21L U103 ( .A(n40), .B(n41), .S(n44), .Z(n39) );
  IVP U104 ( .A(n46), .Z(n45) );
  ND2 U105 ( .A(n108), .B(B[14]), .Z(n107) );
  AN2P U106 ( .A(n106), .B(n22), .Z(n108) );
  EN U107 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  EN U108 ( .A(n7), .B(n49), .Z(SUM[3]) );
  ND2 U109 ( .A(n58), .B(n48), .Z(n7) );
  ND2 U110 ( .A(A[3]), .B(B[3]), .Z(n48) );
  IV U111 ( .A(n47), .Z(n58) );
  MUX21L U112 ( .A(n43), .B(n44), .S(n45), .Z(n42) );
  IV U113 ( .A(n43), .Z(n57) );
  ND2 U114 ( .A(A[6]), .B(B[6]), .Z(n36) );
  MUX21L U115 ( .A(n35), .B(n36), .S(n37), .Z(n34) );
  IV U116 ( .A(n35), .Z(n55) );
  ND2 U117 ( .A(A[4]), .B(B[4]), .Z(n44) );
  ND2 U118 ( .A(A[5]), .B(B[5]), .Z(n41) );
  ND2 U119 ( .A(A[7]), .B(B[7]), .Z(n33) );
endmodule


module prime_DW01_add_78 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n18, n19, n20, n21, n24,
         n25, n26, n29, n30, n31, n32, n33, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n51, n52, n54, n55, n56,
         \A[0] , n103, n104, n105, n106, n107, n108;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  MUX21LP U1 ( .A(n10), .B(n11), .S(n36), .Z(CO) );
  NR2 U4 ( .A(n24), .B(n107), .Z(n12) );
  NR2 U5 ( .A(n25), .B(n107), .Z(n13) );
  NR2 U10 ( .A(n20), .B(n19), .Z(n18) );
  NR2 U19 ( .A(A[8]), .B(B[8]), .Z(n24) );
  MUX21LP U38 ( .A(n38), .B(n37), .S(n45), .Z(n36) );
  FA1A U59 ( .A(n49), .B(A[2]), .CI(B[2]), .CO(n48), .S(SUM[2]) );
  OR2P U68 ( .A(A[6]), .B(B[6]), .Z(n103) );
  MUX21L U69 ( .A(n31), .B(n32), .S(n35), .Z(n30) );
  ND2P U70 ( .A(A[6]), .B(B[6]), .Z(n35) );
  IVA U71 ( .A(n103), .Z(n104) );
  MUX21L U72 ( .A(n31), .B(n32), .S(n105), .Z(n29) );
  NR2P U73 ( .A(A[7]), .B(B[7]), .Z(n31) );
  NR2P U74 ( .A(A[6]), .B(B[6]), .Z(n105) );
  ND2P U75 ( .A(A[4]), .B(B[4]), .Z(n43) );
  EOP U76 ( .A(n36), .B(n5), .Z(SUM[6]) );
  IV U77 ( .A(n55), .Z(n106) );
  IV U78 ( .A(n31), .Z(n52) );
  IV U79 ( .A(n24), .Z(n51) );
  IV U80 ( .A(n42), .Z(n55) );
  NR2P U81 ( .A(A[3]), .B(B[3]), .Z(n46) );
  IV U82 ( .A(n45), .Z(n44) );
  IV U83 ( .A(B[13]), .Z(n19) );
  OR2 U84 ( .A(A[1]), .B(B[1]), .Z(n49) );
  ND2 U85 ( .A(n51), .B(n25), .Z(n3) );
  ND2 U86 ( .A(n52), .B(n32), .Z(n4) );
  ND2 U87 ( .A(A[8]), .B(B[8]), .Z(n25) );
  EN U88 ( .A(n41), .B(n6), .Z(SUM[5]) );
  ND2 U89 ( .A(n54), .B(n40), .Z(n6) );
  EN U90 ( .A(n26), .B(n3), .Z(SUM[8]) );
  EN U91 ( .A(n33), .B(n4), .Z(SUM[7]) );
  IV U92 ( .A(n39), .Z(n54) );
  ND2 U93 ( .A(n56), .B(n47), .Z(n8) );
  MUX21L U94 ( .A(n13), .B(n12), .S(n30), .Z(n11) );
  EO U95 ( .A(n7), .B(n44), .Z(SUM[4]) );
  ND2 U96 ( .A(n55), .B(n43), .Z(n7) );
  ND2 U97 ( .A(n103), .B(n35), .Z(n5) );
  MUX21H U98 ( .A(n29), .B(n30), .S(n36), .Z(n26) );
  AN2P U99 ( .A(B[10]), .B(B[9]), .Z(n21) );
  MUX21L U100 ( .A(n39), .B(n40), .S(n43), .Z(n38) );
  ND2 U101 ( .A(B[11]), .B(B[12]), .Z(n20) );
  ND2 U102 ( .A(n108), .B(B[14]), .Z(n107) );
  AN2P U103 ( .A(n18), .B(n21), .Z(n108) );
  EN U104 ( .A(n8), .B(n48), .Z(SUM[3]) );
  MUX21LP U105 ( .A(n47), .B(n46), .S(n48), .Z(n45) );
  EN U106 ( .A(A[1]), .B(B[1]), .Z(SUM[1]) );
  ND2 U107 ( .A(A[3]), .B(B[3]), .Z(n47) );
  NR2P U108 ( .A(A[5]), .B(B[5]), .Z(n39) );
  IV U109 ( .A(n46), .Z(n56) );
  MUX21L U110 ( .A(n106), .B(n43), .S(n44), .Z(n41) );
  MUX21L U111 ( .A(n39), .B(n40), .S(n42), .Z(n37) );
  NR2P U112 ( .A(A[4]), .B(B[4]), .Z(n42) );
  ND2 U113 ( .A(A[5]), .B(B[5]), .Z(n40) );
  MUX21L U114 ( .A(n104), .B(n35), .S(n36), .Z(n33) );
  MUX21L U115 ( .A(n13), .B(n12), .S(n29), .Z(n10) );
  ND2 U116 ( .A(A[7]), .B(B[7]), .Z(n32) );
endmodule


module prime_DW01_add_76 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1, n5, n6, n11, n15, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n28, n29, n30, n31, n32, \A[0] , n78, n79, n80, n83, n84, n85, n86;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  NR2 U6 ( .A(n78), .B(n11), .Z(n6) );
  NR2 U22 ( .A(A[5]), .B(B[5]), .Z(n21) );
  EOP U24 ( .A(n26), .B(n23), .Z(SUM[4]) );
  MUX21LP U31 ( .A(n30), .B(n31), .S(n1), .Z(n28) );
  FA1AP U44 ( .A(B[2]), .B(A[2]), .CI(n85), .CO(n32), .S(SUM[2]) );
  MUX21LP U45 ( .A(n19), .B(n18), .S(n28), .Z(n15) );
  ND2 U46 ( .A(B[10]), .B(B[9]), .Z(n78) );
  AN2P U47 ( .A(B[8]), .B(B[7]), .Z(n79) );
  ND2P U48 ( .A(A[4]), .B(B[4]), .Z(n25) );
  NR2P U49 ( .A(A[3]), .B(B[3]), .Z(n30) );
  ENP U50 ( .A(A[5]), .B(B[5]), .Z(n20) );
  ENP U51 ( .A(A[4]), .B(B[4]), .Z(n23) );
  NR2P U52 ( .A(A[4]), .B(B[4]), .Z(n24) );
  IVP U53 ( .A(n32), .Z(n1) );
  OR2P U54 ( .A(B[1]), .B(A[1]), .Z(n85) );
  OR2 U55 ( .A(n5), .B(n86), .Z(n80) );
  MUX21L U56 ( .A(n21), .B(n22), .S(n24), .Z(n18) );
  MUX21L U57 ( .A(n21), .B(n22), .S(n25), .Z(n19) );
  EN U58 ( .A(n29), .B(n1), .Z(SUM[3]) );
  EN U59 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  ND2 U60 ( .A(n79), .B(B[6]), .Z(n11) );
  MUX21L U61 ( .A(n83), .B(n84), .S(n28), .Z(SUM[5]) );
  EN U62 ( .A(n20), .B(n25), .Z(n83) );
  EN U63 ( .A(n24), .B(n20), .Z(n84) );
  IV U64 ( .A(n28), .Z(n26) );
  EO U65 ( .A(A[3]), .B(B[3]), .Z(n29) );
  ND2 U66 ( .A(n6), .B(B[11]), .Z(n5) );
  NR2P U67 ( .A(n15), .B(n80), .Z(CO) );
  ND2 U68 ( .A(A[5]), .B(B[5]), .Z(n22) );
  ND2 U69 ( .A(A[3]), .B(B[3]), .Z(n31) );
  IV U70 ( .A(B[12]), .Z(n86) );
endmodule


module prime_DW01_add_97 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n11, n13, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n35, n36, n37, n38, n43, n44, n45, n47,
         n49, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n67, n68, n69, n71, n72, n73, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136;

  AO6P U2 ( .A(n22), .B(n125), .C(n11), .Z(n9) );
  AO6P U6 ( .A(n135), .B(n127), .C(n124), .Z(n13) );
  NR2 U19 ( .A(n32), .B(n27), .Z(n25) );
  NR2 U23 ( .A(A[9]), .B(B[9]), .Z(n27) );
  NR2 U27 ( .A(n134), .B(n32), .Z(n30) );
  NR2 U45 ( .A(A[7]), .B(B[7]), .Z(n43) );
  AO6P U57 ( .A(n52), .B(n60), .C(n53), .Z(n51) );
  NR2 U58 ( .A(n57), .B(n54), .Z(n52) );
  NR2 U68 ( .A(A[4]), .B(B[4]), .Z(n57) );
  FA1A U78 ( .A(n64), .B(A[2]), .CI(B[2]), .CO(n63), .S(SUM[2]) );
  FA1A U79 ( .A(B[1]), .B(A[1]), .CI(n136), .CO(n64), .S(SUM[1]) );
  B3I U87 ( .A(n51), .Z1(n123), .Z2(n122) );
  IV U88 ( .A(n134), .Z(n37) );
  AN2 U89 ( .A(A[11]), .B(B[11]), .Z(n124) );
  AN2 U90 ( .A(n128), .B(n135), .Z(n125) );
  OR2P U91 ( .A(A[6]), .B(B[6]), .Z(n126) );
  AN2 U92 ( .A(A[10]), .B(B[10]), .Z(n127) );
  OR2 U93 ( .A(A[10]), .B(B[10]), .Z(n128) );
  ENP U94 ( .A(n123), .B(n5), .Z(SUM[6]) );
  AO6 U95 ( .A(n123), .B(n37), .C(n132), .Z(n36) );
  AO6 U96 ( .A(n30), .B(n123), .C(n31), .Z(n29) );
  IV U97 ( .A(n72), .Z(n129) );
  NR2P U98 ( .A(A[8]), .B(B[8]), .Z(n32) );
  NR2P U99 ( .A(A[3]), .B(B[3]), .Z(n61) );
  AN2P U100 ( .A(n130), .B(n131), .Z(n54) );
  IVA U101 ( .A(A[5]), .Z(n130) );
  IVDA U102 ( .A(B[5]), .Y(n131) );
  IVDAP U103 ( .A(n38), .Y(n133), .Z(n132) );
  ENP U104 ( .A(n8), .B(n63), .Z(SUM[3]) );
  ND2P U105 ( .A(n126), .B(n69), .Z(n134) );
  IV U106 ( .A(n32), .Z(n68) );
  EOP U107 ( .A(n29), .B(n2), .Z(SUM[9]) );
  EOP U108 ( .A(n36), .B(n3), .Z(SUM[8]) );
  IV U109 ( .A(n49), .Z(n47) );
  AO6P U110 ( .A(n25), .B(n132), .C(n26), .Z(n24) );
  IV U111 ( .A(n60), .Z(n59) );
  ND2 U112 ( .A(n37), .B(n25), .Z(n23) );
  ND2 U113 ( .A(n126), .B(n49), .Z(n5) );
  AO7 U114 ( .A(n43), .B(n49), .C(n44), .Z(n38) );
  IV U115 ( .A(n9), .Z(CO) );
  EO U116 ( .A(n45), .B(n4), .Z(SUM[7]) );
  ND2 U117 ( .A(n69), .B(n44), .Z(n4) );
  AO6 U118 ( .A(n123), .B(n126), .C(n47), .Z(n45) );
  ND2 U119 ( .A(n67), .B(n28), .Z(n2) );
  IV U120 ( .A(n27), .Z(n67) );
  IV U121 ( .A(n43), .Z(n69) );
  IV U122 ( .A(n13), .Z(n11) );
  AO7 U123 ( .A(n122), .B(n23), .C(n24), .Z(n22) );
  ND2 U124 ( .A(A[7]), .B(B[7]), .Z(n44) );
  EO U125 ( .A(n7), .B(n59), .Z(SUM[4]) );
  ND2 U126 ( .A(n72), .B(n58), .Z(n7) );
  ND2 U127 ( .A(A[9]), .B(B[9]), .Z(n28) );
  EN U128 ( .A(n56), .B(n6), .Z(SUM[5]) );
  ND2 U129 ( .A(n71), .B(n55), .Z(n6) );
  AO7 U130 ( .A(n61), .B(n1), .C(n62), .Z(n60) );
  IVP U131 ( .A(n63), .Z(n1) );
  OR2 U132 ( .A(A[11]), .B(B[11]), .Z(n135) );
  ND2 U133 ( .A(n73), .B(n62), .Z(n8) );
  IV U134 ( .A(n61), .Z(n73) );
  OR2 U135 ( .A(B[0]), .B(A[0]), .Z(n136) );
  AO7 U136 ( .A(n59), .B(n129), .C(n58), .Z(n56) );
  IV U137 ( .A(n57), .Z(n72) );
  AO7 U138 ( .A(n54), .B(n58), .C(n55), .Z(n53) );
  IV U139 ( .A(n54), .Z(n71) );
  AO7 U140 ( .A(n133), .B(n32), .C(n35), .Z(n31) );
  ND2 U141 ( .A(n68), .B(n35), .Z(n3) );
  AO7 U142 ( .A(n27), .B(n35), .C(n28), .Z(n26) );
  ND2 U143 ( .A(A[6]), .B(B[6]), .Z(n49) );
  ND2 U144 ( .A(A[8]), .B(B[8]), .Z(n35) );
  EN U145 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  ND2 U146 ( .A(A[5]), .B(B[5]), .Z(n55) );
  ND2 U147 ( .A(A[4]), .B(B[4]), .Z(n58) );
  ND2 U148 ( .A(A[3]), .B(B[3]), .Z(n62) );
endmodule


module prime_DW01_add_95 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n36, n37, n38, n39,
         n40, n41, n44, n45, n46, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n68, n69, n70, n71, n72,
         n73, n74, n123, n124, n125, n126, n127, n128;

  NR2 U10 ( .A(n21), .B(n19), .Z(n17) );
  NR2 U12 ( .A(A[11]), .B(B[11]), .Z(n19) );
  NR2 U14 ( .A(A[10]), .B(B[10]), .Z(n21) );
  NR2 U20 ( .A(n33), .B(n28), .Z(n26) );
  NR2 U28 ( .A(n40), .B(n33), .Z(n31) );
  NR2 U42 ( .A(n49), .B(n44), .Z(n38) );
  NR2 U46 ( .A(A[7]), .B(B[7]), .Z(n44) );
  NR2 U54 ( .A(A[6]), .B(B[6]), .Z(n49) );
  AO6P U58 ( .A(n53), .B(n61), .C(n54), .Z(n52) );
  NR2 U59 ( .A(n58), .B(n55), .Z(n53) );
  NR2 U63 ( .A(A[5]), .B(B[5]), .Z(n55) );
  NR2 U69 ( .A(A[4]), .B(B[4]), .Z(n58) );
  NR2 U77 ( .A(A[3]), .B(B[3]), .Z(n62) );
  FA1A U79 ( .A(n65), .B(A[2]), .CI(B[2]), .CO(n64), .S(SUM[2]) );
  FA1A U80 ( .A(n128), .B(A[1]), .CI(B[1]), .CO(n65), .S(SUM[1]) );
  AN2 U88 ( .A(n18), .B(n127), .Z(n123) );
  AN2 U89 ( .A(n17), .B(n127), .Z(n124) );
  AN2P U90 ( .A(n125), .B(n126), .Z(n28) );
  IV U91 ( .A(A[9]), .Z(n125) );
  IVDA U92 ( .A(B[9]), .Y(n126) );
  ENP U93 ( .A(n8), .B(n64), .Z(SUM[3]) );
  AO7P U94 ( .A(n52), .B(n24), .C(n25), .Z(n23) );
  AO6P U95 ( .A(n26), .B(n39), .C(n27), .Z(n25) );
  IV U96 ( .A(n39), .Z(n41) );
  IV U97 ( .A(n38), .Z(n40) );
  IV U98 ( .A(n50), .Z(n48) );
  IV U99 ( .A(n9), .Z(CO) );
  AO6P U100 ( .A(n23), .B(n124), .C(n123), .Z(n9) );
  IV U101 ( .A(n61), .Z(n60) );
  AO7 U102 ( .A(n44), .B(n50), .C(n45), .Z(n39) );
  AO7 U103 ( .A(n41), .B(n33), .C(n36), .Z(n32) );
  EO U104 ( .A(n37), .B(n3), .Z(SUM[8]) );
  ND2 U105 ( .A(n69), .B(n36), .Z(n3) );
  AO6 U106 ( .A(n51), .B(n38), .C(n39), .Z(n37) );
  IVDA U107 ( .A(n33), .Y(n69) );
  EO U108 ( .A(n46), .B(n4), .Z(SUM[7]) );
  ND2 U109 ( .A(n70), .B(n45), .Z(n4) );
  AO6 U110 ( .A(n51), .B(n71), .C(n48), .Z(n46) );
  IVDA U111 ( .A(n44), .Y(n70) );
  EO U112 ( .A(n30), .B(n2), .Z(SUM[9]) );
  ND2 U113 ( .A(n68), .B(n29), .Z(n2) );
  AO6 U114 ( .A(n51), .B(n31), .C(n32), .Z(n30) );
  ND2 U115 ( .A(A[9]), .B(B[9]), .Z(n29) );
  IV U116 ( .A(n49), .Z(n71) );
  ND2 U117 ( .A(n71), .B(n50), .Z(n5) );
  ND2 U118 ( .A(n26), .B(n38), .Z(n24) );
  ND2 U119 ( .A(A[6]), .B(B[6]), .Z(n50) );
  ND2 U120 ( .A(A[8]), .B(B[8]), .Z(n36) );
  ND2 U121 ( .A(A[7]), .B(B[7]), .Z(n45) );
  IV U122 ( .A(n52), .Z(n51) );
  AN2P U123 ( .A(B[13]), .B(B[12]), .Z(n127) );
  AO7 U124 ( .A(n19), .B(n22), .C(n20), .Z(n18) );
  ND2 U125 ( .A(A[11]), .B(B[11]), .Z(n20) );
  ND2 U126 ( .A(A[10]), .B(B[10]), .Z(n22) );
  EN U127 ( .A(n57), .B(n6), .Z(SUM[5]) );
  EN U128 ( .A(n51), .B(n5), .Z(SUM[6]) );
  ND2 U129 ( .A(n72), .B(n56), .Z(n6) );
  EO U130 ( .A(n7), .B(n60), .Z(SUM[4]) );
  ND2 U131 ( .A(n73), .B(n59), .Z(n7) );
  AO7 U132 ( .A(n62), .B(n1), .C(n63), .Z(n61) );
  IVP U133 ( .A(n64), .Z(n1) );
  ND2 U134 ( .A(n74), .B(n63), .Z(n8) );
  IV U135 ( .A(n62), .Z(n74) );
  OR2 U136 ( .A(B[0]), .B(A[0]), .Z(n128) );
  EN U137 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AO7 U138 ( .A(n28), .B(n36), .C(n29), .Z(n27) );
  IV U139 ( .A(n28), .Z(n68) );
  AO7 U140 ( .A(n60), .B(n58), .C(n59), .Z(n57) );
  IV U141 ( .A(n58), .Z(n73) );
  AO7 U142 ( .A(n55), .B(n59), .C(n56), .Z(n54) );
  IV U143 ( .A(n55), .Z(n72) );
  ND2 U144 ( .A(A[5]), .B(B[5]), .Z(n56) );
  NR2P U145 ( .A(A[8]), .B(B[8]), .Z(n33) );
  ND2 U146 ( .A(A[4]), .B(B[4]), .Z(n59) );
  ND2 U147 ( .A(A[3]), .B(B[3]), .Z(n63) );
endmodule


module prime_DW01_add_98 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n36,
         n37, n38, n39, n40, n41, n44, n45, n46, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n68, n69,
         n70, n71, n72, n73, n74, n123, n124, n125, n126, n127, n128;

  NR2 U7 ( .A(n16), .B(n15), .Z(n14) );
  NR2 U10 ( .A(n21), .B(n19), .Z(n17) );
  NR2 U12 ( .A(A[11]), .B(B[11]), .Z(n19) );
  NR2 U14 ( .A(A[10]), .B(B[10]), .Z(n21) );
  AO7P U17 ( .A(n52), .B(n24), .C(n25), .Z(n23) );
  AO6P U19 ( .A(n26), .B(n39), .C(n27), .Z(n25) );
  NR2 U20 ( .A(n33), .B(n28), .Z(n26) );
  NR2 U24 ( .A(A[9]), .B(B[9]), .Z(n28) );
  NR2 U28 ( .A(n40), .B(n33), .Z(n31) );
  NR2 U42 ( .A(n49), .B(n44), .Z(n38) );
  NR2 U46 ( .A(A[7]), .B(B[7]), .Z(n44) );
  NR2 U54 ( .A(A[6]), .B(B[6]), .Z(n49) );
  NR2 U59 ( .A(n58), .B(n55), .Z(n53) );
  NR2 U69 ( .A(A[4]), .B(B[4]), .Z(n58) );
  ENP U71 ( .A(n8), .B(n64), .Z(SUM[3]) );
  FA1A U79 ( .A(n65), .B(A[2]), .CI(B[2]), .CO(n64), .S(SUM[2]) );
  FA1A U80 ( .A(B[1]), .B(A[1]), .CI(n128), .CO(n65), .S(SUM[1]) );
  AO6 U88 ( .A(n53), .B(n61), .C(n54), .Z(n52) );
  AN2 U89 ( .A(n18), .B(n14), .Z(n123) );
  AO7 U90 ( .A(n1), .B(n62), .C(n63), .Z(n61) );
  IVA U91 ( .A(n61), .Z(n60) );
  AN2 U92 ( .A(n17), .B(n14), .Z(n124) );
  NR2 U93 ( .A(A[3]), .B(B[3]), .Z(n62) );
  NR2P U94 ( .A(A[8]), .B(B[8]), .Z(n33) );
  AO7P U95 ( .A(n125), .B(n60), .C(n126), .Z(n51) );
  IV U96 ( .A(n53), .Z(n125) );
  IV U97 ( .A(n54), .Z(n126) );
  AO7P U98 ( .A(n44), .B(n50), .C(n45), .Z(n39) );
  IVA U99 ( .A(n39), .Z(n41) );
  EOP U100 ( .A(n37), .B(n3), .Z(SUM[8]) );
  EOP U101 ( .A(n46), .B(n4), .Z(SUM[7]) );
  IV U102 ( .A(n73), .Z(n127) );
  ENP U103 ( .A(n51), .B(n5), .Z(SUM[6]) );
  NR2P U104 ( .A(A[5]), .B(B[5]), .Z(n55) );
  AO6P U105 ( .A(n23), .B(n124), .C(n123), .Z(n9) );
  IVA U106 ( .A(n38), .Z(n40) );
  IV U107 ( .A(n50), .Z(n48) );
  IV U108 ( .A(n9), .Z(CO) );
  AO7 U109 ( .A(n28), .B(n36), .C(n29), .Z(n27) );
  EO U110 ( .A(n30), .B(n2), .Z(SUM[9]) );
  ND2 U111 ( .A(n68), .B(n29), .Z(n2) );
  AO6 U112 ( .A(n51), .B(n31), .C(n32), .Z(n30) );
  ND2 U113 ( .A(n69), .B(n36), .Z(n3) );
  AO6 U114 ( .A(n51), .B(n38), .C(n39), .Z(n37) );
  ND2 U115 ( .A(n71), .B(n50), .Z(n5) );
  IV U116 ( .A(n49), .Z(n71) );
  IV U117 ( .A(n28), .Z(n68) );
  ND2 U118 ( .A(n26), .B(n38), .Z(n24) );
  ND2 U119 ( .A(n70), .B(n45), .Z(n4) );
  AO6 U120 ( .A(n51), .B(n71), .C(n48), .Z(n46) );
  ND2 U121 ( .A(A[6]), .B(B[6]), .Z(n50) );
  ND2 U122 ( .A(A[8]), .B(B[8]), .Z(n36) );
  AO7 U123 ( .A(n19), .B(n22), .C(n20), .Z(n18) );
  ND2 U124 ( .A(A[11]), .B(B[11]), .Z(n20) );
  ND2 U125 ( .A(A[10]), .B(B[10]), .Z(n22) );
  ND2 U126 ( .A(A[9]), .B(B[9]), .Z(n29) );
  IV U127 ( .A(n44), .Z(n70) );
  ND2 U128 ( .A(A[7]), .B(B[7]), .Z(n45) );
  EO U129 ( .A(n7), .B(n60), .Z(SUM[4]) );
  ND2 U130 ( .A(n73), .B(n59), .Z(n7) );
  EN U131 ( .A(n57), .B(n6), .Z(SUM[5]) );
  ND2 U132 ( .A(n72), .B(n56), .Z(n6) );
  IVDA U133 ( .A(B[14]), .Y(n15) );
  ND2 U134 ( .A(B[12]), .B(B[13]), .Z(n16) );
  IVP U135 ( .A(n64), .Z(n1) );
  ND2 U136 ( .A(n74), .B(n63), .Z(n8) );
  IV U137 ( .A(n62), .Z(n74) );
  OR2 U138 ( .A(B[0]), .B(A[0]), .Z(n128) );
  EN U139 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AO7 U140 ( .A(n41), .B(n33), .C(n36), .Z(n32) );
  IV U141 ( .A(n33), .Z(n69) );
  AO7 U142 ( .A(n60), .B(n127), .C(n59), .Z(n57) );
  IV U143 ( .A(n58), .Z(n73) );
  AO7 U144 ( .A(n55), .B(n59), .C(n56), .Z(n54) );
  IV U145 ( .A(n55), .Z(n72) );
  ND2 U146 ( .A(A[5]), .B(B[5]), .Z(n56) );
  ND2 U147 ( .A(A[4]), .B(B[4]), .Z(n59) );
  ND2 U148 ( .A(A[3]), .B(B[3]), .Z(n63) );
endmodule


module prime_DW01_add_82 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n17, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n47, n48, n50, n52, \A[0] , n98,
         n99, n100, n101, n102, n103, n104, n105, n106;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  MUX21LP U1 ( .A(n9), .B(n10), .S(n32), .Z(CO) );
  MUX21LP U3 ( .A(n12), .B(n11), .S(n26), .Z(n10) );
  NR2 U5 ( .A(n21), .B(n104), .Z(n12) );
  NR2 U16 ( .A(A[8]), .B(B[8]), .Z(n20) );
  MUX21LP U23 ( .A(n27), .B(n28), .S(n31), .Z(n26) );
  MUX21LP U35 ( .A(n34), .B(n33), .S(n41), .Z(n32) );
  FA1AP U64 ( .A(B[2]), .B(A[2]), .CI(n106), .CO(n44), .S(SUM[2]) );
  IVDA U65 ( .A(n31), .Z(n100) );
  OR2 U66 ( .A(A[4]), .B(B[4]), .Z(n98) );
  MUX21L U67 ( .A(n34), .B(n33), .S(n41), .Z(n99) );
  MUX21LP U68 ( .A(n35), .B(n36), .S(n38), .Z(n33) );
  MUX21LP U69 ( .A(n35), .B(n36), .S(n39), .Z(n34) );
  OR2P U70 ( .A(A[6]), .B(B[6]), .Z(n101) );
  EOP U71 ( .A(n99), .B(n4), .Z(SUM[6]) );
  NR2P U72 ( .A(n20), .B(n104), .Z(n11) );
  ND2P U73 ( .A(A[7]), .B(B[7]), .Z(n28) );
  IV U74 ( .A(n35), .Z(n50) );
  MUX21L U75 ( .A(n12), .B(n11), .S(n25), .Z(n9) );
  MUX21LP U76 ( .A(n27), .B(n28), .S(n30), .Z(n25) );
  IVA U77 ( .A(n25), .Z(n23) );
  NR2P U78 ( .A(A[4]), .B(B[4]), .Z(n38) );
  ND2P U79 ( .A(A[6]), .B(B[6]), .Z(n31) );
  IVA U80 ( .A(n101), .Z(n102) );
  ND2P U81 ( .A(A[4]), .B(B[4]), .Z(n39) );
  NR2 U82 ( .A(A[4]), .B(B[4]), .Z(n103) );
  IV U83 ( .A(n26), .Z(n24) );
  NR2P U84 ( .A(A[7]), .B(B[7]), .Z(n27) );
  NR2P U85 ( .A(A[5]), .B(B[5]), .Z(n35) );
  NR2P U86 ( .A(A[3]), .B(B[3]), .Z(n42) );
  IV U87 ( .A(n41), .Z(n40) );
  OR2P U88 ( .A(B[1]), .B(A[1]), .Z(n106) );
  EN U89 ( .A(n37), .B(n5), .Z(SUM[5]) );
  ND2 U90 ( .A(n98), .B(n39), .Z(n6) );
  EO U91 ( .A(n6), .B(n40), .Z(SUM[4]) );
  MUX21L U92 ( .A(n103), .B(n39), .S(n40), .Z(n37) );
  EN U93 ( .A(n22), .B(n2), .Z(SUM[8]) );
  ND2 U94 ( .A(n47), .B(n21), .Z(n2) );
  MUX21L U95 ( .A(n23), .B(n24), .S(n32), .Z(n22) );
  IV U96 ( .A(n20), .Z(n47) );
  EN U97 ( .A(n29), .B(n3), .Z(SUM[7]) );
  ND2 U98 ( .A(n48), .B(n28), .Z(n3) );
  MUX21L U99 ( .A(n102), .B(n100), .S(n99), .Z(n29) );
  IV U100 ( .A(n27), .Z(n48) );
  ND2 U101 ( .A(n50), .B(n36), .Z(n5) );
  ND2 U102 ( .A(n101), .B(n31), .Z(n4) );
  ND2 U103 ( .A(A[8]), .B(B[8]), .Z(n21) );
  AN2P U104 ( .A(B[10]), .B(B[9]), .Z(n17) );
  MUX21LP U105 ( .A(n43), .B(n42), .S(n44), .Z(n41) );
  EN U106 ( .A(n7), .B(n44), .Z(SUM[3]) );
  ND2 U107 ( .A(n52), .B(n43), .Z(n7) );
  IV U108 ( .A(n42), .Z(n52) );
  ND2 U109 ( .A(n105), .B(B[12]), .Z(n104) );
  AN2P U110 ( .A(n17), .B(B[11]), .Z(n105) );
  EN U111 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  ND2 U112 ( .A(A[3]), .B(B[3]), .Z(n43) );
  ND2 U113 ( .A(A[5]), .B(B[5]), .Z(n36) );
  NR2P U114 ( .A(A[6]), .B(B[6]), .Z(n30) );
endmodule


module prime_DW01_add_79 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n13, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n35, n36, n37,
         n38, n39, n40, n43, n44, n45, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n67, n68, n70, \A[0] ,
         \A[1] , n117, n118, n119, n120, n121, n122, n123, n124, n125, n126;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];

  NR2 U10 ( .A(n20), .B(n18), .Z(n16) );
  NR2 U28 ( .A(n39), .B(n121), .Z(n30) );
  NR2 U42 ( .A(n48), .B(n43), .Z(n37) );
  NR2 U54 ( .A(A[6]), .B(B[6]), .Z(n48) );
  AO6P U58 ( .A(n52), .B(n60), .C(n53), .Z(n51) );
  NR2 U59 ( .A(n57), .B(n54), .Z(n52) );
  NR2 U79 ( .A(B[2]), .B(A[2]), .Z(n63) );
  IVDA U84 ( .A(n57), .Y(n117), .Z(n118) );
  NR2P U85 ( .A(A[4]), .B(B[4]), .Z(n57) );
  ND2P U86 ( .A(A[4]), .B(B[4]), .Z(n58) );
  AO7 U87 ( .A(n18), .B(n21), .C(n19), .Z(n17) );
  AN2 U88 ( .A(n17), .B(n13), .Z(n119) );
  IVDA U89 ( .A(n32), .Y(n120), .Z(n121) );
  AN2 U90 ( .A(n16), .B(n13), .Z(n122) );
  NR2P U91 ( .A(n32), .B(n123), .Z(n25) );
  NR2 U92 ( .A(A[9]), .B(B[9]), .Z(n123) );
  NR2 U93 ( .A(A[9]), .B(B[9]), .Z(n27) );
  EOP U94 ( .A(n29), .B(n1), .Z(SUM[9]) );
  EOP U95 ( .A(n36), .B(n2), .Z(SUM[8]) );
  ND2P U96 ( .A(A[8]), .B(B[8]), .Z(n35) );
  AO7P U97 ( .A(n54), .B(n58), .C(n55), .Z(n53) );
  EOP U98 ( .A(n7), .B(n63), .Z(SUM[3]) );
  OR2 U99 ( .A(A[7]), .B(B[7]), .Z(n125) );
  OR2 U100 ( .A(A[9]), .B(B[9]), .Z(n126) );
  IV U101 ( .A(n38), .Z(n40) );
  AO7P U102 ( .A(n61), .B(n63), .C(n62), .Z(n60) );
  NR2P U103 ( .A(A[3]), .B(B[3]), .Z(n61) );
  NR2P U104 ( .A(A[11]), .B(B[11]), .Z(n18) );
  IVP U105 ( .A(n8), .Z(CO) );
  AO7P U106 ( .A(n43), .B(n49), .C(n44), .Z(n38) );
  ND2 U107 ( .A(A[10]), .B(B[10]), .Z(n21) );
  NR2 U108 ( .A(A[10]), .B(B[10]), .Z(n20) );
  AO6 U109 ( .A(n25), .B(n38), .C(n26), .Z(n24) );
  AO6 U110 ( .A(n22), .B(n122), .C(n119), .Z(n8) );
  IV U111 ( .A(n60), .Z(n59) );
  EOP U112 ( .A(n45), .B(n3), .Z(SUM[7]) );
  ND2 U113 ( .A(n120), .B(n35), .Z(n2) );
  AO7 U114 ( .A(n40), .B(n121), .C(n35), .Z(n31) );
  IV U115 ( .A(n51), .Z(n50) );
  AO7 U116 ( .A(n51), .B(n23), .C(n24), .Z(n22) );
  ND2 U117 ( .A(n126), .B(n28), .Z(n1) );
  AO6 U118 ( .A(n50), .B(n30), .C(n31), .Z(n29) );
  AO6 U119 ( .A(n50), .B(n67), .C(n47), .Z(n45) );
  IVDA U120 ( .A(n49), .Y(n47), .Z(n124) );
  IV U121 ( .A(n48), .Z(n67) );
  ND2 U122 ( .A(n67), .B(n124), .Z(n4) );
  ND2 U123 ( .A(n125), .B(n44), .Z(n3) );
  ND2 U124 ( .A(n70), .B(n62), .Z(n7) );
  ND2 U125 ( .A(A[7]), .B(B[7]), .Z(n44) );
  ND2 U126 ( .A(A[9]), .B(B[9]), .Z(n28) );
  EN U127 ( .A(n56), .B(n5), .Z(SUM[5]) );
  ND2 U128 ( .A(n68), .B(n55), .Z(n5) );
  IV U129 ( .A(n54), .Z(n68) );
  ND2 U130 ( .A(n117), .B(n58), .Z(n6) );
  AN2P U131 ( .A(B[12]), .B(B[13]), .Z(n13) );
  EO U132 ( .A(n6), .B(n59), .Z(SUM[4]) );
  EN U133 ( .A(n50), .B(n4), .Z(SUM[6]) );
  EN U134 ( .A(B[2]), .B(A[2]), .Z(SUM[2]) );
  AO6 U135 ( .A(n50), .B(n37), .C(n38), .Z(n36) );
  IV U136 ( .A(n37), .Z(n39) );
  ND2 U137 ( .A(n25), .B(n37), .Z(n23) );
  AO7 U138 ( .A(n27), .B(n35), .C(n28), .Z(n26) );
  IV U139 ( .A(n61), .Z(n70) );
  ND2 U140 ( .A(A[11]), .B(B[11]), .Z(n19) );
  NR2P U141 ( .A(A[5]), .B(B[5]), .Z(n54) );
  AO7 U142 ( .A(n59), .B(n118), .C(n58), .Z(n56) );
  ND2 U143 ( .A(A[5]), .B(B[5]), .Z(n55) );
  NR2P U144 ( .A(A[8]), .B(B[8]), .Z(n32) );
  ND2 U145 ( .A(A[6]), .B(B[6]), .Z(n49) );
  ND2 U146 ( .A(A[3]), .B(B[3]), .Z(n62) );
  NR2P U147 ( .A(A[7]), .B(B[7]), .Z(n43) );
endmodule


module prime_DW01_add_77 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n10, n11, n13, n14, n15, n16, n18, n60,
         n61;
  assign n14 = B[2];

  NR2 U12 ( .A(n60), .B(n13), .Z(n11) );
  ENP U14 ( .A(n15), .B(n16), .Z(SUM[2]) );
  ND2 U27 ( .A(B[9]), .B(B[8]), .Z(n4) );
  IV U28 ( .A(B[1]), .Z(n61) );
  ND2P U29 ( .A(n7), .B(B[5]), .Z(n6) );
  B4I U30 ( .A(n1), .Z(CO) );
  IV U31 ( .A(n14), .Z(n15) );
  AN2 U32 ( .A(B[7]), .B(B[6]), .Z(n7) );
  ND2 U33 ( .A(n11), .B(B[4]), .Z(n10) );
  ND2 U34 ( .A(n14), .B(n16), .Z(n13) );
  EO U35 ( .A(n61), .B(n18), .Z(SUM[1]) );
  EN U36 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  NR2P U37 ( .A(n6), .B(n10), .Z(n5) );
  NR2P U38 ( .A(n18), .B(n61), .Z(n16) );
  NR2P U39 ( .A(B[0]), .B(A[0]), .Z(n18) );
  ND2P U40 ( .A(n2), .B(n5), .Z(n1) );
  ND2P U41 ( .A(B[10]), .B(B[11]), .Z(n3) );
  NR2P U42 ( .A(n3), .B(n4), .Z(n2) );
  IV U43 ( .A(B[3]), .Z(n60) );
endmodule


module prime_DW01_add_56 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , \A[1] , n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];

  ND2 U36 ( .A(n88), .B(n89), .Z(n80) );
  IVAP U37 ( .A(n70), .Z(CO) );
  B2I U38 ( .A(B[3]), .Z2(n67) );
  IVDAP U39 ( .A(B[4]), .Y(n68), .Z(n69) );
  NR2 U40 ( .A(n92), .B(n93), .Z(n83) );
  ND4P U41 ( .A(n83), .B(n84), .C(n86), .D(n85), .Z(n70) );
  EOP U42 ( .A(A[5]), .B(B[5]), .Z(n74) );
  B3I U43 ( .A(n80), .Z1(n72), .Z2(n71) );
  IVP U44 ( .A(n77), .Z(n73) );
  NR2 U45 ( .A(n76), .B(A[4]), .Z(n75) );
  OR2P U46 ( .A(B[2]), .B(n73), .Z(n82) );
  IVA U47 ( .A(n68), .Z(n76) );
  ND2P U48 ( .A(n69), .B(A[4]), .Z(n81) );
  EO U49 ( .A(n81), .B(n74), .Z(n78) );
  ND2 U50 ( .A(n75), .B(n87), .Z(n86) );
  EO U51 ( .A(n77), .B(B[2]), .Z(SUM[2]) );
  EO U52 ( .A(n75), .B(n74), .Z(n79) );
  ND2 U53 ( .A(B[7]), .B(B[12]), .Z(n93) );
  ND2 U54 ( .A(B[8]), .B(B[11]), .Z(n91) );
  ND2 U55 ( .A(B[6]), .B(B[9]), .Z(n92) );
  ND3P U56 ( .A(n87), .B(n72), .C(n81), .Z(n85) );
  ND2 U57 ( .A(A[3]), .B(n67), .Z(n89) );
  EO3 U58 ( .A(A[3]), .B(n67), .C(n82), .Z(SUM[3]) );
  MUX21L U59 ( .A(n78), .B(n79), .S(n71), .Z(SUM[5]) );
  EO3 U60 ( .A(n69), .B(A[4]), .C(n71), .Z(SUM[4]) );
  AO7 U61 ( .A(A[5]), .B(B[5]), .C(B[10]), .Z(n90) );
  ND2 U62 ( .A(A[5]), .B(B[5]), .Z(n87) );
  IVA U63 ( .A(A[2]), .Z(n77) );
  AO7P U64 ( .A(A[3]), .B(n67), .C(n82), .Z(n88) );
  NR2P U65 ( .A(n90), .B(n91), .Z(n84) );
endmodule


module prime_DW01_add_46 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74;

  EO U30 ( .A(n68), .B(B[0]), .Z(SUM[0]) );
  ND3 U31 ( .A(B[9]), .B(B[8]), .C(B[7]), .Z(n73) );
  IVDAP U32 ( .A(B[2]), .Y(n61), .Z(n62) );
  ENP U33 ( .A(n65), .B(n62), .Z(n67) );
  AO3P U34 ( .A(B[0]), .B(A[0]), .C(B[1]), .D(B[2]), .Z(n71) );
  OR2P U35 ( .A(B[0]), .B(A[0]), .Z(n63) );
  IV U36 ( .A(B[1]), .Z(n64) );
  IVA U37 ( .A(n64), .Z(n65) );
  IVDA U38 ( .A(n63), .Z(n66) );
  EO U39 ( .A(n63), .B(n65), .Z(SUM[1]) );
  MUX21L U40 ( .A(n61), .B(n67), .S(n66), .Z(SUM[2]) );
  AN2P U41 ( .A(n69), .B(n70), .Z(CO) );
  NR2P U42 ( .A(n71), .B(n72), .Z(n70) );
  ND3P U43 ( .A(B[10]), .B(B[4]), .C(B[3]), .Z(n72) );
  IVAP U44 ( .A(A[0]), .Z(n68) );
  NR2P U45 ( .A(n73), .B(n74), .Z(n69) );
  ND2P U46 ( .A(B[6]), .B(B[5]), .Z(n74) );
endmodule


module prime_DW01_add_147 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n5, n8, n12, n13, n14, n15, n16, n17, n18, n19, n21, n22, n25, n26,
         n27, n28, n32, n35, n39, n85, n86, n87, n88, n89, n91, n92, n95, n96,
         n97;

  NR2 U23 ( .A(A[4]), .B(B[4]), .Z(n21) );
  MUX21LP U28 ( .A(n27), .B(n28), .S(n95), .Z(n25) );
  MUX21L U54 ( .A(n18), .B(n19), .S(n22), .Z(n16) );
  OR2 U55 ( .A(B[1]), .B(A[1]), .Z(n85) );
  OR2P U56 ( .A(B[0]), .B(A[0]), .Z(n86) );
  AN2P U57 ( .A(B[2]), .B(A[2]), .Z(n87) );
  AN2P U58 ( .A(B[1]), .B(A[1]), .Z(n88) );
  OR2 U59 ( .A(n5), .B(n97), .Z(n89) );
  MUX21H U60 ( .A(n14), .B(n13), .S(n25), .Z(SUM[5]) );
  AN2P U61 ( .A(B[8]), .B(B[9]), .Z(n91) );
  NR2P U62 ( .A(n12), .B(n89), .Z(CO) );
  EOP U63 ( .A(A[3]), .B(B[3]), .Z(n26) );
  ENP U64 ( .A(A[5]), .B(B[5]), .Z(n17) );
  NR2 U65 ( .A(A[5]), .B(B[5]), .Z(n18) );
  MUX21LP U66 ( .A(n92), .B(n87), .S(n35), .Z(n95) );
  OR2 U67 ( .A(B[2]), .B(A[2]), .Z(n92) );
  EN U68 ( .A(n26), .B(n95), .Z(SUM[3]) );
  EO U69 ( .A(n39), .B(n86), .Z(SUM[1]) );
  EN U70 ( .A(n35), .B(n32), .Z(SUM[2]) );
  MUX21L U71 ( .A(n16), .B(n15), .S(n25), .Z(n12) );
  EO U72 ( .A(n17), .B(n22), .Z(n14) );
  EN U73 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  MUX21L U74 ( .A(n88), .B(n85), .S(n86), .Z(n35) );
  MUX21L U75 ( .A(n18), .B(n19), .S(n21), .Z(n15) );
  EO U76 ( .A(n21), .B(n17), .Z(n13) );
  EO U77 ( .A(B[2]), .B(A[2]), .Z(n32) );
  EO U78 ( .A(B[1]), .B(A[1]), .Z(n39) );
  EO U79 ( .A(n25), .B(n96), .Z(SUM[4]) );
  EO U80 ( .A(A[4]), .B(B[4]), .Z(n96) );
  NR2 U81 ( .A(A[3]), .B(B[3]), .Z(n27) );
  ND2 U82 ( .A(A[4]), .B(B[4]), .Z(n22) );
  AN2P U83 ( .A(B[6]), .B(B[7]), .Z(n8) );
  ND2 U84 ( .A(n8), .B(n91), .Z(n5) );
  ND2 U85 ( .A(A[3]), .B(B[3]), .Z(n28) );
  ND2 U86 ( .A(A[5]), .B(B[5]), .Z(n19) );
  IV U87 ( .A(B[10]), .Z(n97) );
endmodule


module prime_DW01_add_114 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n18, n19, n20, n21, n22,
         n23, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n48, n49, n51, n53, \A[0] ,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  MUX21LP U1 ( .A(n10), .B(n11), .S(n33), .Z(CO) );
  NR2 U10 ( .A(n20), .B(n19), .Z(n18) );
  ND2P U14 ( .A(n48), .B(n22), .Z(n3) );
  NR2 U16 ( .A(A[8]), .B(B[8]), .Z(n21) );
  ENP U34 ( .A(n6), .B(n38), .Z(SUM[5]) );
  EOP U42 ( .A(n7), .B(n41), .Z(SUM[4]) );
  ENP U48 ( .A(n8), .B(n45), .Z(SUM[3]) );
  FA1A U56 ( .A(n46), .B(A[2]), .CI(B[2]), .CO(n45), .S(SUM[2]) );
  IVDA U65 ( .A(n34), .Z(n98) );
  IVDA U66 ( .A(n35), .Z(n99) );
  MUX21L U67 ( .A(n36), .B(n37), .S(n40), .Z(n35) );
  MUX21L U68 ( .A(n36), .B(n37), .S(n39), .Z(n34) );
  MUX21LP U69 ( .A(n35), .B(n34), .S(n42), .Z(n33) );
  NR2P U70 ( .A(A[3]), .B(B[3]), .Z(n43) );
  OR2 U71 ( .A(A[4]), .B(B[4]), .Z(n100) );
  ND2P U72 ( .A(A[4]), .B(B[4]), .Z(n40) );
  OR2 U73 ( .A(A[6]), .B(B[6]), .Z(n101) );
  MUX21L U74 ( .A(n28), .B(n29), .S(n32), .Z(n27) );
  NR2P U75 ( .A(A[7]), .B(B[7]), .Z(n28) );
  IVA U76 ( .A(n100), .Z(n102) );
  NR2P U77 ( .A(n21), .B(n105), .Z(n12) );
  NR2P U78 ( .A(n22), .B(n105), .Z(n13) );
  MUX21LP U79 ( .A(n99), .B(n98), .S(n42), .Z(n103) );
  EOP U80 ( .A(n103), .B(n5), .Z(SUM[6]) );
  ND2P U81 ( .A(A[6]), .B(B[6]), .Z(n32) );
  IVA U82 ( .A(n101), .Z(n104) );
  MUX21L U83 ( .A(n28), .B(n29), .S(n31), .Z(n26) );
  IV U84 ( .A(n42), .Z(n41) );
  EN U85 ( .A(n23), .B(n3), .Z(SUM[8]) );
  MUX21L U86 ( .A(n13), .B(n12), .S(n27), .Z(n11) );
  MUX21H U87 ( .A(n26), .B(n27), .S(n103), .Z(n23) );
  IV U88 ( .A(n21), .Z(n48) );
  ND2 U89 ( .A(n51), .B(n37), .Z(n6) );
  IV U90 ( .A(n36), .Z(n51) );
  ND2 U91 ( .A(n106), .B(B[13]), .Z(n105) );
  AN2P U92 ( .A(n18), .B(B[12]), .Z(n106) );
  ND2 U93 ( .A(A[8]), .B(B[8]), .Z(n22) );
  EN U94 ( .A(n30), .B(n4), .Z(SUM[7]) );
  ND2 U95 ( .A(n49), .B(n29), .Z(n4) );
  IV U96 ( .A(n28), .Z(n49) );
  IVP U97 ( .A(B[11]), .Z(n19) );
  ND2 U98 ( .A(A[3]), .B(B[3]), .Z(n44) );
  MUX21LP U99 ( .A(n44), .B(n43), .S(n45), .Z(n42) );
  ND2 U100 ( .A(n53), .B(n44), .Z(n8) );
  EN U101 ( .A(A[1]), .B(B[1]), .Z(SUM[1]) );
  IVP U102 ( .A(A[1]), .Z(n107) );
  IV U103 ( .A(B[1]), .Z(n108) );
  ND2P U104 ( .A(n107), .B(n108), .Z(n46) );
  ND2 U105 ( .A(A[5]), .B(B[5]), .Z(n37) );
  IV U106 ( .A(n43), .Z(n53) );
  ND2 U107 ( .A(B[10]), .B(B[9]), .Z(n20) );
  ND2 U108 ( .A(n101), .B(n32), .Z(n5) );
  ND2 U109 ( .A(n100), .B(n40), .Z(n7) );
  MUX21L U110 ( .A(n13), .B(n12), .S(n26), .Z(n10) );
  ND2 U111 ( .A(A[7]), .B(B[7]), .Z(n29) );
  NR2P U112 ( .A(A[5]), .B(B[5]), .Z(n36) );
  MUX21L U113 ( .A(n102), .B(n40), .S(n41), .Z(n38) );
  NR2P U114 ( .A(A[4]), .B(B[4]), .Z(n39) );
  MUX21L U115 ( .A(n104), .B(n32), .S(n103), .Z(n30) );
  NR2P U116 ( .A(A[6]), .B(B[6]), .Z(n31) );
endmodule


module prime_DW01_add_104 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n12, n13, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n35, n36, n37, n38, n39, n40, n43, n44, n45,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n66, n68, n69, n70, n71, n72, \A[0] , n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  AO6P U6 ( .A(n126), .B(n118), .C(n124), .Z(n13) );
  EOP U15 ( .A(n29), .B(n2), .Z(SUM[9]) );
  AO7P U16 ( .A(n51), .B(n23), .C(n24), .Z(n22) );
  AO6P U18 ( .A(n25), .B(n38), .C(n26), .Z(n24) );
  NR2 U27 ( .A(n39), .B(n121), .Z(n30) );
  AO6P U57 ( .A(n52), .B(n60), .C(n53), .Z(n51) );
  NR2 U68 ( .A(A[4]), .B(B[4]), .Z(n57) );
  NR2 U76 ( .A(A[3]), .B(B[3]), .Z(n61) );
  FA1A U78 ( .A(B[2]), .B(A[2]), .CI(n127), .CO(n63), .S(SUM[2]) );
  OR2P U86 ( .A(A[8]), .B(B[8]), .Z(n125) );
  IVAP U87 ( .A(n125), .Z(n121) );
  AN2 U88 ( .A(A[10]), .B(B[10]), .Z(n118) );
  OR2 U89 ( .A(A[10]), .B(B[10]), .Z(n119) );
  OR2P U90 ( .A(A[11]), .B(B[11]), .Z(n126) );
  AO7P U91 ( .A(n120), .B(n12), .C(n13), .Z(CO) );
  IV U92 ( .A(n22), .Z(n120) );
  NR2P U93 ( .A(n57), .B(n54), .Z(n52) );
  AO7 U94 ( .A(n54), .B(n58), .C(n55), .Z(n53) );
  NR2P U95 ( .A(A[5]), .B(B[5]), .Z(n54) );
  NR2P U96 ( .A(n43), .B(n48), .Z(n37) );
  NR2 U97 ( .A(A[6]), .B(B[6]), .Z(n48) );
  NR2P U98 ( .A(n27), .B(n121), .Z(n25) );
  AO7P U99 ( .A(n61), .B(n1), .C(n62), .Z(n60) );
  NR2 U100 ( .A(n27), .B(n121), .Z(n122) );
  NR2P U101 ( .A(A[9]), .B(B[9]), .Z(n27) );
  NR2P U102 ( .A(A[7]), .B(B[7]), .Z(n43) );
  IV U103 ( .A(n40), .Z(n123) );
  AO7 U104 ( .A(n43), .B(n49), .C(n44), .Z(n38) );
  IV U105 ( .A(n38), .Z(n40) );
  IV U106 ( .A(n37), .Z(n39) );
  AO6P U107 ( .A(n30), .B(n50), .C(n31), .Z(n29) );
  IV U108 ( .A(n60), .Z(n59) );
  AN2 U109 ( .A(A[11]), .B(B[11]), .Z(n124) );
  AO6 U110 ( .A(n50), .B(n69), .C(n47), .Z(n45) );
  IV U111 ( .A(n48), .Z(n69) );
  IV U112 ( .A(n51), .Z(n50) );
  EO U113 ( .A(n45), .B(n4), .Z(SUM[7]) );
  EO U114 ( .A(n36), .B(n3), .Z(SUM[8]) );
  AO6 U115 ( .A(n50), .B(n37), .C(n123), .Z(n36) );
  EN U116 ( .A(n56), .B(n6), .Z(SUM[5]) );
  ND2 U117 ( .A(n70), .B(n55), .Z(n6) );
  ND2 U118 ( .A(n125), .B(n35), .Z(n3) );
  EO U119 ( .A(n7), .B(n59), .Z(SUM[4]) );
  ND2 U120 ( .A(n71), .B(n58), .Z(n7) );
  ND2 U121 ( .A(n66), .B(n28), .Z(n2) );
  EN U122 ( .A(n50), .B(n5), .Z(SUM[6]) );
  ND2 U123 ( .A(n68), .B(n44), .Z(n4) );
  IVP U124 ( .A(n63), .Z(n1) );
  EN U125 ( .A(n8), .B(n63), .Z(SUM[3]) );
  ND2 U126 ( .A(n72), .B(n62), .Z(n8) );
  ND2 U127 ( .A(n119), .B(n126), .Z(n12) );
  OR2 U128 ( .A(B[1]), .B(A[1]), .Z(n127) );
  EN U129 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  ND2 U130 ( .A(n69), .B(n49), .Z(n5) );
  IV U131 ( .A(n49), .Z(n47) );
  IV U132 ( .A(n61), .Z(n72) );
  ND2 U133 ( .A(A[8]), .B(B[8]), .Z(n35) );
  AO7 U134 ( .A(n59), .B(n57), .C(n58), .Z(n56) );
  IV U135 ( .A(n57), .Z(n71) );
  AO7 U136 ( .A(n27), .B(n35), .C(n28), .Z(n26) );
  IV U137 ( .A(n27), .Z(n66) );
  IV U138 ( .A(n43), .Z(n68) );
  ND2 U139 ( .A(A[6]), .B(B[6]), .Z(n49) );
  IV U140 ( .A(n54), .Z(n70) );
  ND2 U141 ( .A(A[7]), .B(B[7]), .Z(n44) );
  ND2 U142 ( .A(A[5]), .B(B[5]), .Z(n55) );
  ND2 U143 ( .A(A[3]), .B(B[3]), .Z(n62) );
  AO7 U144 ( .A(n40), .B(n121), .C(n35), .Z(n31) );
  ND2 U145 ( .A(n122), .B(n37), .Z(n23) );
  ND2 U146 ( .A(A[9]), .B(B[9]), .Z(n28) );
  ND2 U147 ( .A(A[4]), .B(B[4]), .Z(n58) );
endmodule


module prime_DW01_add_116 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n18, n19, n20, n21, n22,
         n23, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n41, n42, n43, n44, n45, n46, n48, n49, n50, n51, n52, n53, n98,
         n99, n100, n101, n102, n103;

  NR2 U4 ( .A(n21), .B(n101), .Z(n12) );
  NR2 U5 ( .A(n22), .B(n101), .Z(n13) );
  NR2 U10 ( .A(n20), .B(n19), .Z(n18) );
  NR2 U16 ( .A(A[8]), .B(B[8]), .Z(n21) );
  ENP U18 ( .A(n30), .B(n4), .Z(SUM[7]) );
  EOP U28 ( .A(n33), .B(n5), .Z(SUM[6]) );
  ENP U34 ( .A(n6), .B(n38), .Z(SUM[5]) );
  MUX21LP U35 ( .A(n35), .B(n34), .S(n42), .Z(n33) );
  EOP U42 ( .A(n7), .B(n41), .Z(SUM[4]) );
  ENP U48 ( .A(n8), .B(n45), .Z(SUM[3]) );
  NR2 U54 ( .A(A[3]), .B(B[3]), .Z(n43) );
  FA1A U57 ( .A(n103), .B(A[1]), .CI(B[1]), .CO(n46), .S(SUM[1]) );
  ND2P U65 ( .A(A[4]), .B(B[4]), .Z(n98) );
  IVP U66 ( .A(n52), .Z(n99) );
  FA1AP U67 ( .A(B[2]), .B(A[2]), .CI(n46), .CO(n45), .S(SUM[2]) );
  IVA U68 ( .A(n50), .Z(n100) );
  MUX21LP U69 ( .A(n10), .B(n11), .S(n33), .Z(CO) );
  MUX21L U70 ( .A(n36), .B(n37), .S(n98), .Z(n35) );
  MUX21L U71 ( .A(n36), .B(n37), .S(n39), .Z(n34) );
  NR2P U72 ( .A(A[5]), .B(B[5]), .Z(n36) );
  NR2P U73 ( .A(A[4]), .B(B[4]), .Z(n39) );
  ENP U74 ( .A(n23), .B(n3), .Z(SUM[8]) );
  IV U75 ( .A(n36), .Z(n51) );
  IV U76 ( .A(n39), .Z(n52) );
  IV U77 ( .A(n42), .Z(n41) );
  IV U78 ( .A(B[11]), .Z(n19) );
  MUX21L U79 ( .A(n28), .B(n29), .S(n31), .Z(n26) );
  MUX21L U80 ( .A(n28), .B(n29), .S(n32), .Z(n27) );
  ND2 U81 ( .A(n48), .B(n22), .Z(n3) );
  IV U82 ( .A(n21), .Z(n48) );
  ND2 U83 ( .A(n49), .B(n29), .Z(n4) );
  IV U84 ( .A(n28), .Z(n49) );
  ND2 U85 ( .A(n50), .B(n32), .Z(n5) );
  IV U86 ( .A(n31), .Z(n50) );
  MUX21L U87 ( .A(n13), .B(n12), .S(n27), .Z(n11) );
  MUX21L U88 ( .A(n13), .B(n12), .S(n26), .Z(n10) );
  MUX21H U89 ( .A(n26), .B(n27), .S(n33), .Z(n23) );
  ND2 U90 ( .A(A[8]), .B(B[8]), .Z(n22) );
  MUX21L U91 ( .A(n100), .B(n32), .S(n33), .Z(n30) );
  ND2 U92 ( .A(n52), .B(n98), .Z(n7) );
  ND2 U93 ( .A(n51), .B(n37), .Z(n6) );
  MUX21L U94 ( .A(n99), .B(n98), .S(n41), .Z(n38) );
  EN U95 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  ND2 U96 ( .A(A[3]), .B(B[3]), .Z(n44) );
  ND2 U97 ( .A(B[9]), .B(B[10]), .Z(n20) );
  ND2 U98 ( .A(n102), .B(B[13]), .Z(n101) );
  AN2P U99 ( .A(n18), .B(B[12]), .Z(n102) );
  MUX21LP U100 ( .A(n44), .B(n43), .S(n45), .Z(n42) );
  ND2 U101 ( .A(n53), .B(n44), .Z(n8) );
  IV U102 ( .A(n43), .Z(n53) );
  OR2 U103 ( .A(B[0]), .B(A[0]), .Z(n103) );
  ND2 U104 ( .A(A[5]), .B(B[5]), .Z(n37) );
  NR2P U105 ( .A(A[7]), .B(B[7]), .Z(n28) );
  NR2P U106 ( .A(A[6]), .B(B[6]), .Z(n31) );
  ND2 U107 ( .A(A[7]), .B(B[7]), .Z(n29) );
  ND2 U108 ( .A(A[6]), .B(B[6]), .Z(n32) );
endmodule


module prime_DW01_add_126 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n48, n49, n50, n51,
         n52, n98, n99, n100, n101, n102, n103, n104, n105;

  NR2 U4 ( .A(n20), .B(n103), .Z(n11) );
  NR2 U5 ( .A(n21), .B(n103), .Z(n12) );
  NR2 U10 ( .A(n19), .B(n18), .Z(n17) );
  ENP U13 ( .A(n22), .B(n2), .Z(SUM[8]) );
  ND2P U14 ( .A(n48), .B(n21), .Z(n2) );
  NR2 U16 ( .A(A[8]), .B(B[8]), .Z(n20) );
  ENP U18 ( .A(n29), .B(n3), .Z(SUM[7]) );
  ENP U34 ( .A(n5), .B(n37), .Z(SUM[5]) );
  MUX21LP U35 ( .A(n34), .B(n33), .S(n41), .Z(n32) );
  EOP U42 ( .A(n6), .B(n40), .Z(SUM[4]) );
  ENP U48 ( .A(n7), .B(n44), .Z(SUM[3]) );
  NR2 U54 ( .A(A[3]), .B(B[3]), .Z(n42) );
  FA1A U57 ( .A(B[1]), .B(A[1]), .CI(n105), .CO(n45), .S(SUM[1]) );
  B2I U65 ( .A(n33), .Z2(n98) );
  MUX21L U66 ( .A(n35), .B(n36), .S(n38), .Z(n33) );
  ND2P U67 ( .A(A[4]), .B(B[4]), .Z(n39) );
  MUX21LP U68 ( .A(n34), .B(n98), .S(n41), .Z(n99) );
  IVA U69 ( .A(n52), .Z(n100) );
  IV U70 ( .A(n38), .Z(n52) );
  MUX21L U71 ( .A(n9), .B(n10), .S(n32), .Z(CO) );
  IVA U72 ( .A(n50), .Z(n101) );
  MUX21L U73 ( .A(n27), .B(n28), .S(n30), .Z(n25) );
  ND2P U74 ( .A(A[6]), .B(B[6]), .Z(n31) );
  NR2P U75 ( .A(A[5]), .B(B[5]), .Z(n35) );
  IV U76 ( .A(n25), .Z(n23) );
  MUX21LP U77 ( .A(n27), .B(n28), .S(n31), .Z(n26) );
  IV U78 ( .A(n30), .Z(n50) );
  IV U79 ( .A(n43), .Z(n102) );
  NR2P U80 ( .A(A[4]), .B(B[4]), .Z(n38) );
  IV U81 ( .A(n41), .Z(n40) );
  OR2P U82 ( .A(B[0]), .B(A[0]), .Z(n105) );
  IVP U83 ( .A(n26), .Z(n24) );
  MUX21L U84 ( .A(n12), .B(n11), .S(n26), .Z(n10) );
  MUX21L U85 ( .A(n12), .B(n11), .S(n25), .Z(n9) );
  MUX21L U86 ( .A(n23), .B(n24), .S(n99), .Z(n22) );
  IV U87 ( .A(n20), .Z(n48) );
  ND2 U88 ( .A(n52), .B(n39), .Z(n6) );
  ND2 U89 ( .A(n49), .B(n28), .Z(n3) );
  MUX21L U90 ( .A(n101), .B(n31), .S(n99), .Z(n29) );
  IV U91 ( .A(n27), .Z(n49) );
  MUX21L U92 ( .A(n100), .B(n39), .S(n40), .Z(n37) );
  ND2 U93 ( .A(n50), .B(n31), .Z(n4) );
  OR2 U94 ( .A(n42), .B(n102), .Z(n7) );
  ND2 U95 ( .A(n51), .B(n36), .Z(n5) );
  IVP U96 ( .A(n35), .Z(n51) );
  ND2 U97 ( .A(n104), .B(B[13]), .Z(n103) );
  AN2P U98 ( .A(n17), .B(B[12]), .Z(n104) );
  EO U99 ( .A(n32), .B(n4), .Z(SUM[6]) );
  EN U100 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  MUX21L U101 ( .A(n35), .B(n36), .S(n39), .Z(n34) );
  ND2 U102 ( .A(A[3]), .B(B[3]), .Z(n43) );
  ND2 U103 ( .A(A[8]), .B(B[8]), .Z(n21) );
  IV U104 ( .A(B[11]), .Z(n18) );
  ND2 U105 ( .A(B[10]), .B(B[9]), .Z(n19) );
  MUX21LP U106 ( .A(n43), .B(n42), .S(n44), .Z(n41) );
  FA1A U107 ( .A(B[2]), .B(A[2]), .CI(n45), .CO(n44), .S(SUM[2]) );
  ND2 U108 ( .A(A[5]), .B(B[5]), .Z(n36) );
  NR2P U109 ( .A(A[7]), .B(B[7]), .Z(n27) );
  ND2 U110 ( .A(A[7]), .B(B[7]), .Z(n28) );
  NR2P U111 ( .A(A[6]), .B(B[6]), .Z(n30) );
endmodule


module prime_DW01_add_121 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n14, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n39, n40, n41,
         n42, n46, n47, n48, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n70, n72, n75, n76, n123,
         n125, n126, n127, n128, n129, n130, n131, n132;

  NR2 U12 ( .A(A[11]), .B(B[11]), .Z(n19) );
  NR2 U14 ( .A(A[10]), .B(B[10]), .Z(n21) );
  MUX21LP U17 ( .A(n24), .B(n25), .S(n54), .Z(n23) );
  NR2 U24 ( .A(A[9]), .B(B[9]), .Z(n28) );
  NR2 U36 ( .A(A[8]), .B(B[8]), .Z(n33) );
  FA1A U81 ( .A(B[2]), .B(A[2]), .CI(n67), .CO(n66), .S(SUM[2]) );
  FA1A U82 ( .A(n132), .B(A[1]), .CI(B[1]), .CO(n67), .S(SUM[1]) );
  MUX21H U90 ( .A(n127), .B(n125), .S(n23), .Z(CO) );
  AN2P U91 ( .A(n17), .B(n14), .Z(n125) );
  B2I U92 ( .A(n33), .Z1(n123), .Z2(n126) );
  AN2 U93 ( .A(n18), .B(n14), .Z(n127) );
  IVA U94 ( .A(n128), .Z(n57) );
  IVAP U95 ( .A(n54), .Z(n53) );
  NR2P U96 ( .A(A[3]), .B(B[3]), .Z(n64) );
  OR2P U97 ( .A(A[5]), .B(B[5]), .Z(n128) );
  IVDA U98 ( .A(n61), .Z(n129) );
  IV U99 ( .A(n75), .Z(n130) );
  OR2 U100 ( .A(A[6]), .B(B[6]), .Z(n131) );
  NR2 U101 ( .A(A[6]), .B(B[6]), .Z(n51) );
  IVAP U102 ( .A(n40), .Z(n42) );
  NR2P U103 ( .A(A[4]), .B(B[4]), .Z(n60) );
  MUX21LP U104 ( .A(n46), .B(n47), .S(n52), .Z(n41) );
  NR2P U105 ( .A(A[7]), .B(B[7]), .Z(n46) );
  MUX21LP U106 ( .A(n46), .B(n47), .S(n51), .Z(n40) );
  MUX21LP U107 ( .A(n28), .B(n29), .S(n126), .Z(n26) );
  MUX21L U108 ( .A(n28), .B(n29), .S(n34), .Z(n27) );
  ND2 U109 ( .A(n76), .B(n65), .Z(n8) );
  IV U110 ( .A(n46), .Z(n72) );
  EOP U111 ( .A(n39), .B(n3), .Z(SUM[8]) );
  MUX21L U112 ( .A(n34), .B(n126), .S(n41), .Z(n32) );
  IV U113 ( .A(n64), .Z(n76) );
  MUX21LP U114 ( .A(n56), .B(n55), .S(n63), .Z(n54) );
  MUX21LP U115 ( .A(n65), .B(n64), .S(n66), .Z(n63) );
  MUX21L U116 ( .A(n27), .B(n26), .S(n40), .Z(n24) );
  MUX21L U117 ( .A(n27), .B(n26), .S(n41), .Z(n25) );
  MUX21L U118 ( .A(n50), .B(n131), .S(n53), .Z(n48) );
  IVDA U119 ( .A(n52), .Y(n50) );
  MUX21L U120 ( .A(n41), .B(n40), .S(n53), .Z(n39) );
  ND2 U121 ( .A(n131), .B(n52), .Z(n5) );
  ND2 U122 ( .A(n72), .B(n47), .Z(n4) );
  EO U123 ( .A(n30), .B(n2), .Z(SUM[9]) );
  EO U124 ( .A(n48), .B(n4), .Z(SUM[7]) );
  EN U125 ( .A(n53), .B(n5), .Z(SUM[6]) );
  EN U126 ( .A(n59), .B(n6), .Z(SUM[5]) );
  MUX21L U127 ( .A(n32), .B(n31), .S(n53), .Z(n30) );
  MUX21L U128 ( .A(n126), .B(n34), .S(n42), .Z(n31) );
  ND2 U129 ( .A(n70), .B(n29), .Z(n2) );
  IV U130 ( .A(n28), .Z(n70) );
  EO U131 ( .A(n7), .B(n62), .Z(SUM[4]) );
  ND2 U132 ( .A(n128), .B(n58), .Z(n6) );
  ND2 U133 ( .A(n123), .B(n34), .Z(n3) );
  ND2 U134 ( .A(n75), .B(n61), .Z(n7) );
  MUX21L U135 ( .A(n57), .B(n58), .S(n61), .Z(n56) );
  MUX21L U136 ( .A(n57), .B(n58), .S(n60), .Z(n55) );
  MUX21L U137 ( .A(n19), .B(n20), .S(n21), .Z(n17) );
  IVP U138 ( .A(n63), .Z(n62) );
  MUX21L U139 ( .A(n19), .B(n20), .S(n22), .Z(n18) );
  ND2 U140 ( .A(A[10]), .B(B[10]), .Z(n22) );
  ND2 U141 ( .A(A[11]), .B(B[11]), .Z(n20) );
  AN2P U142 ( .A(B[13]), .B(B[12]), .Z(n14) );
  EN U143 ( .A(n8), .B(n66), .Z(SUM[3]) );
  EN U144 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  OR2 U145 ( .A(B[0]), .B(A[0]), .Z(n132) );
  MUX21L U146 ( .A(n130), .B(n129), .S(n62), .Z(n59) );
  IV U147 ( .A(n60), .Z(n75) );
  ND2 U148 ( .A(A[8]), .B(B[8]), .Z(n34) );
  ND2 U149 ( .A(A[6]), .B(B[6]), .Z(n52) );
  ND2 U150 ( .A(A[3]), .B(B[3]), .Z(n65) );
  ND2 U151 ( .A(A[7]), .B(B[7]), .Z(n47) );
  ND2 U152 ( .A(A[9]), .B(B[9]), .Z(n29) );
  ND2 U153 ( .A(A[5]), .B(B[5]), .Z(n58) );
  ND2 U154 ( .A(A[4]), .B(B[4]), .Z(n61) );
endmodule


module prime_DW01_add_123 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n39, n40, n41, n46,
         n47, n48, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n70, n73, n74, n76, n123, n124, n125,
         n126, n127, n128, n129, n131, n132;

  NR2 U12 ( .A(A[11]), .B(B[11]), .Z(n19) );
  NR2 U14 ( .A(A[10]), .B(B[10]), .Z(n21) );
  NR2 U36 ( .A(A[8]), .B(B[8]), .Z(n33) );
  FA1A U81 ( .A(n67), .B(A[2]), .CI(B[2]), .CO(n66), .S(SUM[2]) );
  FA1A U82 ( .A(n132), .B(A[1]), .CI(B[1]), .CO(n67), .S(SUM[1]) );
  IVA U90 ( .A(n129), .Z(n60) );
  B2I U91 ( .A(n33), .Z1(n123), .Z2(n124) );
  AN2 U92 ( .A(n17), .B(B[12]), .Z(n125) );
  NR2P U93 ( .A(A[9]), .B(B[9]), .Z(n28) );
  NR2P U94 ( .A(A[6]), .B(B[6]), .Z(n51) );
  MUX21L U95 ( .A(n58), .B(n57), .S(n129), .Z(n55) );
  NR2 U96 ( .A(A[7]), .B(B[7]), .Z(n46) );
  OR2P U97 ( .A(A[7]), .B(B[7]), .Z(n126) );
  AN2P U98 ( .A(A[7]), .B(B[7]), .Z(n127) );
  MUX21LP U99 ( .A(n126), .B(n127), .S(n51), .Z(n128) );
  B4I U100 ( .A(n128), .Z(n40) );
  NR2P U101 ( .A(A[3]), .B(B[3]), .Z(n64) );
  ENP U102 ( .A(n53), .B(n5), .Z(SUM[6]) );
  MUX21LP U103 ( .A(n28), .B(n29), .S(n124), .Z(n26) );
  MUX21LP U104 ( .A(n27), .B(n26), .S(n41), .Z(n25) );
  OR2P U105 ( .A(A[4]), .B(B[4]), .Z(n129) );
  MUX21LP U106 ( .A(n46), .B(n47), .S(n52), .Z(n41) );
  MUX21LP U107 ( .A(n57), .B(n58), .S(n61), .Z(n56) );
  NR2P U108 ( .A(A[5]), .B(B[5]), .Z(n57) );
  IVAP U109 ( .A(n54), .Z(n53) );
  MUX21LP U110 ( .A(n19), .B(n20), .S(n21), .Z(n17) );
  EOP U111 ( .A(n39), .B(n3), .Z(SUM[8]) );
  MUX21H U112 ( .A(n131), .B(n125), .S(n23), .Z(CO) );
  MUX21L U113 ( .A(n34), .B(n124), .S(n41), .Z(n32) );
  MUX21LP U114 ( .A(n56), .B(n55), .S(n63), .Z(n54) );
  AN2 U115 ( .A(n18), .B(B[12]), .Z(n131) );
  IV U116 ( .A(n64), .Z(n76) );
  MUX21LP U117 ( .A(n65), .B(n64), .S(n66), .Z(n63) );
  MUX21L U118 ( .A(n41), .B(n40), .S(n53), .Z(n39) );
  EO U119 ( .A(n30), .B(n2), .Z(SUM[9]) );
  ND2 U120 ( .A(n70), .B(n29), .Z(n2) );
  EO U121 ( .A(n48), .B(n4), .Z(SUM[7]) );
  ND2 U122 ( .A(n126), .B(n47), .Z(n4) );
  ND2 U123 ( .A(n123), .B(n34), .Z(n3) );
  ND2 U124 ( .A(n73), .B(n52), .Z(n5) );
  MUX21L U125 ( .A(n24), .B(n25), .S(n54), .Z(n23) );
  MUX21L U126 ( .A(n27), .B(n26), .S(n40), .Z(n24) );
  MUX21L U127 ( .A(n28), .B(n29), .S(n34), .Z(n27) );
  EN U128 ( .A(n59), .B(n6), .Z(SUM[5]) );
  ND2 U129 ( .A(n74), .B(n58), .Z(n6) );
  MUX21L U130 ( .A(n32), .B(n31), .S(n53), .Z(n30) );
  MUX21L U131 ( .A(n124), .B(n34), .S(n128), .Z(n31) );
  MUX21L U132 ( .A(n50), .B(n73), .S(n53), .Z(n48) );
  IV U133 ( .A(n52), .Z(n50) );
  IV U134 ( .A(n51), .Z(n73) );
  IV U135 ( .A(n28), .Z(n70) );
  EO U136 ( .A(n7), .B(n62), .Z(SUM[4]) );
  ND2 U137 ( .A(n129), .B(n61), .Z(n7) );
  IV U138 ( .A(n57), .Z(n74) );
  ND2 U139 ( .A(A[11]), .B(B[11]), .Z(n20) );
  IVP U140 ( .A(n63), .Z(n62) );
  MUX21L U141 ( .A(n19), .B(n20), .S(n22), .Z(n18) );
  ND2 U142 ( .A(A[10]), .B(B[10]), .Z(n22) );
  EN U143 ( .A(n8), .B(n66), .Z(SUM[3]) );
  ND2 U144 ( .A(n76), .B(n65), .Z(n8) );
  EN U145 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  OR2 U146 ( .A(B[0]), .B(A[0]), .Z(n132) );
  MUX21L U147 ( .A(n60), .B(n61), .S(n62), .Z(n59) );
  ND2 U148 ( .A(A[8]), .B(B[8]), .Z(n34) );
  ND2 U149 ( .A(A[6]), .B(B[6]), .Z(n52) );
  ND2 U150 ( .A(A[3]), .B(B[3]), .Z(n65) );
  ND2 U151 ( .A(A[7]), .B(B[7]), .Z(n47) );
  ND2 U152 ( .A(A[9]), .B(B[9]), .Z(n29) );
  ND2 U153 ( .A(A[5]), .B(B[5]), .Z(n58) );
  ND2 U154 ( .A(A[4]), .B(B[4]), .Z(n61) );
endmodule


module prime_DW01_add_141 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n6, n7, n9, n12, n13, n14, n15, n16, n18, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n50, n51, n52, n53,
         n55, n58, n59, n60, n61, n62, n64, n65, n68, n70, n71, n72, n76, n77,
         n78, \B[0] , n129, n130, n131, n133, n134, n135, n136, n137, n139;
  assign n9 = B[11];
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  MUX21LP U2 ( .A(n135), .B(n130), .S(n23), .Z(SUM[12]) );
  NR2 U7 ( .A(n14), .B(n131), .Z(n6) );
  NR2 U8 ( .A(n15), .B(n131), .Z(n7) );
  MUX21LP U13 ( .A(n13), .B(n12), .S(n23), .Z(SUM[11]) );
  EOP U14 ( .A(n21), .B(n16), .Z(n12) );
  EOP U15 ( .A(n16), .B(n22), .Z(n13) );
  NR2 U24 ( .A(A[10]), .B(B[10]), .Z(n21) );
  MUX21LP U27 ( .A(n26), .B(n27), .S(n55), .Z(n23) );
  MUX21LP U39 ( .A(n36), .B(n35), .S(n53), .Z(SUM[8]) );
  EOP U40 ( .A(n40), .B(n37), .Z(n35) );
  EOP U41 ( .A(n41), .B(n37), .Z(n36) );
  MUX21LP U50 ( .A(n47), .B(n48), .S(n51), .Z(n44) );
  MUX21LP U51 ( .A(n47), .B(n48), .S(n52), .Z(n45) );
  NR2 U53 ( .A(A[7]), .B(B[7]), .Z(n47) );
  MUX21LP U63 ( .A(n59), .B(n58), .S(n68), .Z(n55) );
  MUX21LP U67 ( .A(n61), .B(n62), .S(n65), .Z(n59) );
  NR2 U69 ( .A(B[5]), .B(A[5]), .Z(n61) );
  NR2 U73 ( .A(B[4]), .B(A[4]), .Z(n64) );
  MUX21LP U78 ( .A(n70), .B(n71), .S(n72), .Z(n68) );
  NR2 U80 ( .A(B[3]), .B(A[3]), .Z(n70) );
  NR2 U88 ( .A(B[2]), .B(A[2]), .Z(n77) );
  EOP U96 ( .A(B[2]), .B(A[2]), .Z(n76) );
  NR2P U97 ( .A(A[11]), .B(n131), .Z(n129) );
  EOP U98 ( .A(n14), .B(n131), .Z(n130) );
  IVDAP U99 ( .A(n9), .Z(n131) );
  ENP U100 ( .A(A[1]), .B(B[1]), .Z(SUM[1]) );
  EOP U101 ( .A(n51), .B(n46), .Z(n42) );
  MUX21LP U102 ( .A(n7), .B(n6), .S(n23), .Z(SUM[13]) );
  NR2P U103 ( .A(A[6]), .B(B[6]), .Z(n51) );
  ND2 U104 ( .A(A[9]), .B(B[9]), .Z(n34) );
  ENP U105 ( .A(A[9]), .B(B[9]), .Z(n32) );
  NR2 U106 ( .A(A[9]), .B(B[9]), .Z(n33) );
  EOP U107 ( .A(n15), .B(n131), .Z(n135) );
  ND2 U108 ( .A(B[8]), .B(A[8]), .Z(n39) );
  NR2 U109 ( .A(B[8]), .B(A[8]), .Z(n38) );
  EOP U110 ( .A(A[6]), .B(B[6]), .Z(n50) );
  EOP U111 ( .A(B[8]), .B(A[8]), .Z(n37) );
  EOP U112 ( .A(A[10]), .B(B[10]), .Z(n20) );
  EOP U113 ( .A(A[11]), .B(n131), .Z(n16) );
  IV U114 ( .A(n45), .Z(n41) );
  IV U115 ( .A(n44), .Z(n40) );
  OR2P U116 ( .A(A[1]), .B(B[1]), .Z(n136) );
  MUX21L U117 ( .A(n61), .B(n62), .S(n64), .Z(n58) );
  MUX21LP U118 ( .A(n129), .B(n18), .S(n21), .Z(n14) );
  MUX21L U119 ( .A(n31), .B(n30), .S(n45), .Z(n27) );
  MUX21L U120 ( .A(n31), .B(n30), .S(n44), .Z(n26) );
  MUX21L U121 ( .A(n33), .B(n34), .S(n39), .Z(n31) );
  MUX21L U122 ( .A(n133), .B(n134), .S(n68), .Z(SUM[5]) );
  EN U123 ( .A(n60), .B(n65), .Z(n133) );
  EN U124 ( .A(n60), .B(n64), .Z(n134) );
  MUX21L U125 ( .A(n24), .B(n25), .S(n55), .Z(SUM[9]) );
  MUX21L U126 ( .A(n29), .B(n28), .S(n45), .Z(n25) );
  MUX21L U127 ( .A(n29), .B(n28), .S(n44), .Z(n24) );
  EO U128 ( .A(n32), .B(n39), .Z(n29) );
  IV U129 ( .A(n55), .Z(n53) );
  MUX21L U130 ( .A(n33), .B(n34), .S(n38), .Z(n30) );
  EO U131 ( .A(n38), .B(n32), .Z(n28) );
  ND2 U132 ( .A(B[5]), .B(A[5]), .Z(n62) );
  MUX21H U133 ( .A(n78), .B(n77), .S(n136), .Z(n72) );
  ND2 U134 ( .A(B[2]), .B(A[2]), .Z(n78) );
  MUX21L U135 ( .A(n129), .B(n18), .S(n22), .Z(n15) );
  EOP U136 ( .A(n53), .B(n50), .Z(SUM[6]) );
  ND2 U137 ( .A(A[7]), .B(B[7]), .Z(n48) );
  MUX21L U138 ( .A(n43), .B(n42), .S(n53), .Z(SUM[7]) );
  EO U139 ( .A(n46), .B(n52), .Z(n43) );
  EO U140 ( .A(A[7]), .B(B[7]), .Z(n46) );
  EN U141 ( .A(B[5]), .B(A[5]), .Z(n60) );
  EO U142 ( .A(n68), .B(n137), .Z(SUM[4]) );
  EO U143 ( .A(B[4]), .B(A[4]), .Z(n137) );
  EO U144 ( .A(n76), .B(n136), .Z(SUM[2]) );
  EO U145 ( .A(n139), .B(n72), .Z(SUM[3]) );
  EN U146 ( .A(B[3]), .B(A[3]), .Z(n139) );
  ND2 U147 ( .A(B[4]), .B(A[4]), .Z(n65) );
  EOP U148 ( .A(n23), .B(n20), .Z(SUM[10]) );
  ND2 U149 ( .A(A[11]), .B(n131), .Z(n18) );
  ND2 U150 ( .A(A[6]), .B(B[6]), .Z(n52) );
  ND2 U151 ( .A(B[3]), .B(A[3]), .Z(n71) );
  ND2 U152 ( .A(A[10]), .B(B[10]), .Z(n22) );
endmodule


module prime_DW01_add_111 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n31, n32,
         n33, \A[0] , n76, n77;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  NR2 U6 ( .A(n13), .B(n12), .Z(n11) );
  NR2 U9 ( .A(n16), .B(n15), .Z(n14) );
  ENP U12 ( .A(n22), .B(n3), .Z(SUM[5]) );
  AO6P U13 ( .A(n18), .B(n26), .C(n19), .Z(n17) );
  NR2 U14 ( .A(n23), .B(n20), .Z(n18) );
  NR2 U18 ( .A(A[5]), .B(B[5]), .Z(n20) );
  NR2 U24 ( .A(A[4]), .B(B[4]), .Z(n23) );
  ENP U26 ( .A(n5), .B(n29), .Z(SUM[3]) );
  AO7P U28 ( .A(n27), .B(n1), .C(n28), .Z(n26) );
  FA1A U34 ( .A(n77), .B(A[2]), .CI(B[2]), .CO(n29), .S(SUM[2]) );
  IV U42 ( .A(n32), .Z(n76) );
  ND2P U43 ( .A(B[12]), .B(B[11]), .Z(n10) );
  NR2P U44 ( .A(A[3]), .B(B[3]), .Z(n27) );
  NR2P U45 ( .A(n10), .B(n9), .Z(n8) );
  ND2P U46 ( .A(B[14]), .B(B[13]), .Z(n9) );
  IV U47 ( .A(B[6]), .Z(n16) );
  IV U48 ( .A(B[7]), .Z(n15) );
  AO7 U49 ( .A(n20), .B(n24), .C(n21), .Z(n19) );
  ND2 U50 ( .A(n14), .B(B[8]), .Z(n13) );
  ND2 U51 ( .A(B[9]), .B(B[10]), .Z(n12) );
  ND2 U52 ( .A(n31), .B(n21), .Z(n3) );
  IV U53 ( .A(n20), .Z(n31) );
  ND2 U54 ( .A(n32), .B(n24), .Z(n4) );
  IV U55 ( .A(n26), .Z(n25) );
  IV U56 ( .A(n29), .Z(n1) );
  EO U57 ( .A(n25), .B(n4), .Z(SUM[4]) );
  EN U58 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  ND2 U59 ( .A(n33), .B(n28), .Z(n5) );
  IV U60 ( .A(n27), .Z(n33) );
  OR2 U61 ( .A(B[1]), .B(A[1]), .Z(n77) );
  AO7 U62 ( .A(n25), .B(n76), .C(n24), .Z(n22) );
  IV U63 ( .A(n23), .Z(n32) );
  ND2 U64 ( .A(A[5]), .B(B[5]), .Z(n21) );
  ND2 U65 ( .A(A[4]), .B(B[4]), .Z(n24) );
  ND2 U66 ( .A(A[3]), .B(B[3]), .Z(n28) );
  NR2P U67 ( .A(n7), .B(n17), .Z(CO) );
  ND2 U68 ( .A(n8), .B(n11), .Z(n7) );
endmodule


module prime_DW01_add_138 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1, n4, n5, n6, n7, n8, n9, n10, n12, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n25, n26, n27, n28, n29, n30, n77, n78, n79;

  NR2 U1 ( .A(n4), .B(n12), .Z(CO) );
  NR2 U6 ( .A(n10), .B(n9), .Z(n8) );
  MUX21LP U11 ( .A(n16), .B(n15), .S(n25), .Z(n12) );
  NR2 U17 ( .A(A[5]), .B(B[5]), .Z(n18) );
  EOP U19 ( .A(n23), .B(n20), .Z(SUM[4]) );
  NR2 U21 ( .A(A[4]), .B(B[4]), .Z(n21) );
  MUX21LP U26 ( .A(n27), .B(n28), .S(n1), .Z(n25) );
  NR2 U28 ( .A(A[3]), .B(B[3]), .Z(n27) );
  FA1A U31 ( .A(n30), .B(A[2]), .CI(B[2]), .CO(n29), .S(SUM[2]) );
  FA1A U32 ( .A(n79), .B(A[1]), .CI(B[1]), .CO(n30), .S(SUM[1]) );
  NR2P U40 ( .A(n6), .B(n7), .Z(n5) );
  ND2P U41 ( .A(B[13]), .B(B[12]), .Z(n6) );
  ENP U42 ( .A(A[5]), .B(B[5]), .Z(n17) );
  ENP U43 ( .A(A[4]), .B(B[4]), .Z(n20) );
  ND2P U44 ( .A(B[7]), .B(B[6]), .Z(n10) );
  IVAP U45 ( .A(n29), .Z(n1) );
  MUX21L U46 ( .A(n18), .B(n19), .S(n22), .Z(n16) );
  ND2P U47 ( .A(B[11]), .B(B[10]), .Z(n7) );
  ND2 U48 ( .A(B[8]), .B(B[9]), .Z(n9) );
  MUX21L U49 ( .A(n18), .B(n19), .S(n21), .Z(n15) );
  ND2 U50 ( .A(n5), .B(n8), .Z(n4) );
  EN U51 ( .A(n26), .B(n1), .Z(SUM[3]) );
  MUX21L U52 ( .A(n77), .B(n78), .S(n25), .Z(SUM[5]) );
  EN U53 ( .A(n17), .B(n22), .Z(n77) );
  EN U54 ( .A(n21), .B(n17), .Z(n78) );
  IV U55 ( .A(n25), .Z(n23) );
  ND2 U56 ( .A(A[3]), .B(B[3]), .Z(n28) );
  OR2 U57 ( .A(B[0]), .B(A[0]), .Z(n79) );
  EO U58 ( .A(A[3]), .B(B[3]), .Z(n26) );
  EN U59 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  ND2 U60 ( .A(A[5]), .B(B[5]), .Z(n19) );
  ND2 U61 ( .A(A[4]), .B(B[4]), .Z(n22) );
endmodule


module prime_DW01_add_100 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36,
         n37, n40, n41, n42, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n63, n64, n66, n67, \A[0] , \A[1] ,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];

  NR2 U7 ( .A(n17), .B(n15), .Z(n13) );
  NR2 U11 ( .A(A[10]), .B(B[10]), .Z(n17) );
  AO7P U14 ( .A(n48), .B(n20), .C(n21), .Z(n19) );
  AO6P U16 ( .A(n22), .B(n35), .C(n23), .Z(n21) );
  EOP U23 ( .A(n33), .B(n2), .Z(SUM[8]) );
  NR2 U25 ( .A(n36), .B(n121), .Z(n27) );
  EOP U33 ( .A(n42), .B(n3), .Z(SUM[7]) );
  ND2P U52 ( .A(A[6]), .B(B[6]), .Z(n46) );
  AO6P U55 ( .A(n49), .B(n57), .C(n50), .Z(n48) );
  NR2 U56 ( .A(n54), .B(n51), .Z(n49) );
  EOP U62 ( .A(n6), .B(n56), .Z(SUM[4]) );
  NR2 U66 ( .A(A[4]), .B(B[4]), .Z(n54) );
  EOP U68 ( .A(n7), .B(n60), .Z(SUM[3]) );
  AO7P U70 ( .A(n58), .B(n60), .C(n59), .Z(n57) );
  NR2 U76 ( .A(B[2]), .B(A[2]), .Z(n60) );
  NR2P U81 ( .A(n29), .B(n24), .Z(n22) );
  NR2P U82 ( .A(A[11]), .B(B[11]), .Z(n15) );
  AN2 U83 ( .A(n13), .B(B[12]), .Z(n112) );
  NR2 U84 ( .A(A[9]), .B(B[9]), .Z(n113) );
  NR2 U85 ( .A(A[9]), .B(B[9]), .Z(n24) );
  NR2P U86 ( .A(A[7]), .B(B[7]), .Z(n40) );
  B5I U87 ( .A(n114), .Z(CO) );
  AO6P U88 ( .A(n19), .B(n112), .C(n123), .Z(n114) );
  NR2P U89 ( .A(A[8]), .B(B[8]), .Z(n29) );
  ND2 U90 ( .A(A[3]), .B(B[3]), .Z(n59) );
  NR2 U91 ( .A(A[7]), .B(B[7]), .Z(n122) );
  OR2 U92 ( .A(A[8]), .B(B[8]), .Z(n115) );
  OR2 U93 ( .A(A[9]), .B(B[9]), .Z(n116) );
  AO7 U94 ( .A(n113), .B(n32), .C(n25), .Z(n23) );
  ND2P U95 ( .A(A[8]), .B(B[8]), .Z(n32) );
  AO7P U96 ( .A(n40), .B(n46), .C(n41), .Z(n35) );
  ND2 U97 ( .A(A[7]), .B(B[7]), .Z(n41) );
  OR2 U98 ( .A(A[5]), .B(B[5]), .Z(n117) );
  IV U99 ( .A(n66), .Z(n118) );
  B2I U100 ( .A(n32), .Z2(n119) );
  IV U101 ( .A(n37), .Z(n120) );
  IVA U102 ( .A(n115), .Z(n121) );
  AO7P U103 ( .A(n51), .B(n55), .C(n52), .Z(n50) );
  ENP U104 ( .A(n53), .B(n5), .Z(SUM[5]) );
  NR2P U105 ( .A(A[5]), .B(B[5]), .Z(n51) );
  AN2 U106 ( .A(n14), .B(B[12]), .Z(n123) );
  ND2 U107 ( .A(n63), .B(n41), .Z(n3) );
  AO6 U108 ( .A(n47), .B(n64), .C(n44), .Z(n42) );
  EN U109 ( .A(n47), .B(n4), .Z(SUM[6]) );
  ND2 U110 ( .A(n64), .B(n46), .Z(n4) );
  IV U111 ( .A(n45), .Z(n64) );
  ND2 U112 ( .A(n67), .B(n59), .Z(n7) );
  IV U113 ( .A(n58), .Z(n67) );
  EO U114 ( .A(n26), .B(n1), .Z(SUM[9]) );
  ND2 U115 ( .A(n116), .B(n25), .Z(n1) );
  AO6 U116 ( .A(n47), .B(n27), .C(n28), .Z(n26) );
  IV U117 ( .A(n57), .Z(n56) );
  ND2 U118 ( .A(n115), .B(n119), .Z(n2) );
  AO7 U119 ( .A(n15), .B(n18), .C(n16), .Z(n14) );
  ND2 U120 ( .A(A[10]), .B(B[10]), .Z(n18) );
  EN U121 ( .A(B[2]), .B(A[2]), .Z(SUM[2]) );
  IV U122 ( .A(n34), .Z(n36) );
  IV U123 ( .A(n48), .Z(n47) );
  IV U124 ( .A(n46), .Z(n44) );
  IV U125 ( .A(n122), .Z(n63) );
  AO6 U126 ( .A(n47), .B(n34), .C(n120), .Z(n33) );
  IV U127 ( .A(n35), .Z(n37) );
  AO7 U128 ( .A(n37), .B(n121), .C(n119), .Z(n28) );
  IV U129 ( .A(n54), .Z(n66) );
  ND2 U130 ( .A(n66), .B(n55), .Z(n6) );
  ND2 U131 ( .A(n117), .B(n52), .Z(n5) );
  ND2 U132 ( .A(A[11]), .B(B[11]), .Z(n16) );
  ND2 U133 ( .A(n22), .B(n34), .Z(n20) );
  ND2 U134 ( .A(A[9]), .B(B[9]), .Z(n25) );
  ND2 U135 ( .A(A[5]), .B(B[5]), .Z(n52) );
  ND2 U136 ( .A(A[4]), .B(B[4]), .Z(n55) );
  NR2P U137 ( .A(n45), .B(n122), .Z(n34) );
  NR2P U138 ( .A(A[6]), .B(B[6]), .Z(n45) );
  NR2P U139 ( .A(A[3]), .B(B[3]), .Z(n58) );
  AO7 U140 ( .A(n56), .B(n118), .C(n55), .Z(n53) );
endmodule


module prime_DW01_add_149 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n5, n6, n7, n8, n10, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n23, n25, n26, n27, \A[0] , n71, n72, n74, n75, n77, n78;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  NR2 U6 ( .A(n8), .B(n7), .Z(n6) );
  NR2 U17 ( .A(A[5]), .B(B[5]), .Z(n16) );
  MUX21LP U26 ( .A(n25), .B(n26), .S(n1), .Z(n23) );
  OR2 U39 ( .A(n5), .B(n78), .Z(n71) );
  FA1 U40 ( .A(B[2]), .B(A[2]), .CI(n72), .CO(n27), .S(SUM[2]) );
  NR2P U41 ( .A(A[4]), .B(B[4]), .Z(n19) );
  MUX21L U42 ( .A(n14), .B(n13), .S(n23), .Z(n10) );
  ENP U43 ( .A(n19), .B(n15), .Z(n75) );
  ENP U44 ( .A(A[5]), .B(B[5]), .Z(n15) );
  NR2P U45 ( .A(A[3]), .B(B[3]), .Z(n25) );
  IV U46 ( .A(n27), .Z(n1) );
  OR2P U47 ( .A(B[1]), .B(A[1]), .Z(n72) );
  NR2P U48 ( .A(n10), .B(n71), .Z(CO) );
  MUX21L U49 ( .A(n74), .B(n75), .S(n23), .Z(SUM[5]) );
  EN U50 ( .A(n15), .B(n20), .Z(n74) );
  IV U51 ( .A(n23), .Z(n21) );
  EN U52 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  EN U53 ( .A(A[4]), .B(B[4]), .Z(n18) );
  ND2 U54 ( .A(B[8]), .B(B[9]), .Z(n7) );
  EO U55 ( .A(n77), .B(n1), .Z(SUM[3]) );
  EN U56 ( .A(A[3]), .B(B[3]), .Z(n77) );
  ND2 U57 ( .A(B[7]), .B(B[6]), .Z(n8) );
  MUX21L U58 ( .A(n16), .B(n17), .S(n19), .Z(n13) );
  EO U59 ( .A(n21), .B(n18), .Z(SUM[4]) );
  MUX21L U60 ( .A(n16), .B(n17), .S(n20), .Z(n14) );
  ND2 U61 ( .A(n6), .B(B[10]), .Z(n5) );
  ND2 U62 ( .A(A[3]), .B(B[3]), .Z(n26) );
  ND2 U63 ( .A(A[4]), .B(B[4]), .Z(n20) );
  ND2 U64 ( .A(A[5]), .B(B[5]), .Z(n17) );
  IV U65 ( .A(B[11]), .Z(n78) );
endmodule


module prime_DW01_add_134 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n12, n13, n14, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n34, n40, n41,
         n46, n47, n48, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n70, n71, n72, n73, n74, n75, n76,
         n123, n124, n126, n127;

  NR2 U12 ( .A(A[11]), .B(B[11]), .Z(n19) );
  NR2 U14 ( .A(A[10]), .B(B[10]), .Z(n21) );
  NR2 U24 ( .A(A[9]), .B(B[9]), .Z(n28) );
  NR2 U48 ( .A(A[7]), .B(B[7]), .Z(n46) );
  NR2 U56 ( .A(A[6]), .B(B[6]), .Z(n51) );
  NR2 U65 ( .A(A[5]), .B(B[5]), .Z(n57) );
  NR2 U71 ( .A(A[4]), .B(B[4]), .Z(n60) );
  NR2 U79 ( .A(A[3]), .B(B[3]), .Z(n64) );
  FA1A U81 ( .A(B[2]), .B(A[2]), .CI(n67), .CO(n66), .S(SUM[2]) );
  FA1A U82 ( .A(B[1]), .B(A[1]), .CI(n127), .CO(n67), .S(SUM[1]) );
  MUX21L U90 ( .A(n24), .B(n25), .S(n54), .Z(n23) );
  ND2P U91 ( .A(A[8]), .B(B[8]), .Z(n34) );
  IVA U92 ( .A(n71), .Z(n123) );
  NR2 U93 ( .A(A[8]), .B(B[8]), .Z(n124) );
  MUX21L U94 ( .A(n13), .B(n12), .S(n23), .Z(CO) );
  MUX21LP U95 ( .A(n46), .B(n47), .S(n51), .Z(n40) );
  MUX21LP U96 ( .A(n28), .B(n29), .S(n34), .Z(n27) );
  ENP U97 ( .A(n126), .B(n3), .Z(SUM[8]) );
  MUX21H U98 ( .A(n41), .B(n40), .S(n53), .Z(n126) );
  MUX21LP U99 ( .A(n56), .B(n55), .S(n63), .Z(n54) );
  ND2P U100 ( .A(n17), .B(n14), .Z(n12) );
  MUX21LP U101 ( .A(n65), .B(n64), .S(n66), .Z(n63) );
  EN U102 ( .A(n59), .B(n6), .Z(SUM[5]) );
  EO U103 ( .A(n48), .B(n4), .Z(SUM[7]) );
  ND2 U104 ( .A(n72), .B(n47), .Z(n4) );
  MUX21L U105 ( .A(n50), .B(n73), .S(n53), .Z(n48) );
  IV U106 ( .A(n46), .Z(n72) );
  EO U107 ( .A(n7), .B(n62), .Z(SUM[4]) );
  MUX21L U108 ( .A(n46), .B(n47), .S(n52), .Z(n41) );
  MUX21L U109 ( .A(n28), .B(n29), .S(n124), .Z(n26) );
  MUX21L U110 ( .A(n27), .B(n26), .S(n40), .Z(n24) );
  MUX21L U111 ( .A(n27), .B(n26), .S(n41), .Z(n25) );
  IVP U112 ( .A(n54), .Z(n53) );
  EO U113 ( .A(n30), .B(n2), .Z(SUM[9]) );
  ND2 U114 ( .A(n70), .B(n29), .Z(n2) );
  MUX21L U115 ( .A(n32), .B(n31), .S(n53), .Z(n30) );
  IV U116 ( .A(n28), .Z(n70) );
  ND2 U117 ( .A(n71), .B(n34), .Z(n3) );
  IV U118 ( .A(n124), .Z(n71) );
  MUX21L U119 ( .A(n34), .B(n123), .S(n40), .Z(n31) );
  MUX21L U120 ( .A(n34), .B(n123), .S(n41), .Z(n32) );
  EN U121 ( .A(n53), .B(n5), .Z(SUM[6]) );
  ND2 U122 ( .A(n73), .B(n52), .Z(n5) );
  ND2 U123 ( .A(A[11]), .B(B[11]), .Z(n20) );
  IV U124 ( .A(n52), .Z(n50) );
  MUX21L U125 ( .A(n60), .B(n61), .S(n62), .Z(n59) );
  ND2 U126 ( .A(n74), .B(n58), .Z(n6) );
  IV U127 ( .A(n57), .Z(n74) );
  ND2 U128 ( .A(n75), .B(n61), .Z(n7) );
  IV U129 ( .A(n60), .Z(n75) );
  AN2P U130 ( .A(B[12]), .B(B[13]), .Z(n14) );
  MUX21L U131 ( .A(n57), .B(n58), .S(n61), .Z(n56) );
  MUX21L U132 ( .A(n57), .B(n58), .S(n60), .Z(n55) );
  ND2 U133 ( .A(n18), .B(n14), .Z(n13) );
  MUX21L U134 ( .A(n19), .B(n20), .S(n22), .Z(n18) );
  ND2 U135 ( .A(A[10]), .B(B[10]), .Z(n22) );
  MUX21L U136 ( .A(n19), .B(n20), .S(n21), .Z(n17) );
  IVP U137 ( .A(n63), .Z(n62) );
  EN U138 ( .A(n8), .B(n66), .Z(SUM[3]) );
  ND2 U139 ( .A(n76), .B(n65), .Z(n8) );
  IV U140 ( .A(n64), .Z(n76) );
  OR2 U141 ( .A(B[0]), .B(A[0]), .Z(n127) );
  EN U142 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  IV U143 ( .A(n51), .Z(n73) );
  ND2 U144 ( .A(A[6]), .B(B[6]), .Z(n52) );
  ND2 U145 ( .A(A[3]), .B(B[3]), .Z(n65) );
  ND2 U146 ( .A(A[7]), .B(B[7]), .Z(n47) );
  ND2 U147 ( .A(A[9]), .B(B[9]), .Z(n29) );
  ND2 U148 ( .A(A[5]), .B(B[5]), .Z(n58) );
  ND2 U149 ( .A(A[4]), .B(B[4]), .Z(n61) );
endmodule


module prime_DW01_add_133 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n29, n30, n31, n32, n33, n34, n37, n38, n39, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n61, n62, n63, n64, n65, n66, n67, n114, n115, n116,
         n117;

  NR2 U13 ( .A(n26), .B(n21), .Z(n19) );
  NR2 U17 ( .A(A[9]), .B(B[9]), .Z(n21) );
  NR2 U21 ( .A(n33), .B(n26), .Z(n24) );
  NR2 U27 ( .A(A[8]), .B(B[8]), .Z(n26) );
  NR2 U35 ( .A(n42), .B(n37), .Z(n31) );
  NR2 U47 ( .A(A[6]), .B(B[6]), .Z(n42) );
  AO6P U51 ( .A(n46), .B(n54), .C(n47), .Z(n45) );
  NR2 U52 ( .A(n51), .B(n48), .Z(n46) );
  NR2 U56 ( .A(A[5]), .B(B[5]), .Z(n48) );
  NR2 U62 ( .A(A[4]), .B(B[4]), .Z(n51) );
  NR2 U70 ( .A(A[3]), .B(B[3]), .Z(n55) );
  FA1A U72 ( .A(B[2]), .B(A[2]), .CI(n58), .CO(n57), .S(SUM[2]) );
  FA1A U73 ( .A(B[1]), .B(A[1]), .CI(n117), .CO(n58), .S(SUM[1]) );
  OR2 U81 ( .A(A[10]), .B(B[10]), .Z(n114) );
  OR2 U82 ( .A(n116), .B(A[11]), .Z(n115) );
  NR2 U83 ( .A(A[7]), .B(B[7]), .Z(n37) );
  IV U84 ( .A(n45), .Z(n44) );
  IV U85 ( .A(n9), .Z(CO) );
  IV U86 ( .A(n31), .Z(n33) );
  IV U87 ( .A(n54), .Z(n53) );
  AN2 U88 ( .A(A[10]), .B(B[10]), .Z(n116) );
  EO U89 ( .A(n39), .B(n4), .Z(SUM[7]) );
  ND2 U90 ( .A(n63), .B(n38), .Z(n4) );
  AO6 U91 ( .A(n44), .B(n64), .C(n41), .Z(n39) );
  IV U92 ( .A(n37), .Z(n63) );
  EN U93 ( .A(n50), .B(n6), .Z(SUM[5]) );
  ND2 U94 ( .A(n65), .B(n49), .Z(n6) );
  AO7 U95 ( .A(n53), .B(n51), .C(n52), .Z(n50) );
  IV U96 ( .A(n48), .Z(n65) );
  EO U97 ( .A(n7), .B(n53), .Z(SUM[4]) );
  ND2 U98 ( .A(n66), .B(n52), .Z(n7) );
  IV U99 ( .A(n51), .Z(n66) );
  AO7 U100 ( .A(n37), .B(n43), .C(n38), .Z(n32) );
  AO7 U101 ( .A(n48), .B(n52), .C(n49), .Z(n47) );
  AO7 U102 ( .A(n45), .B(n17), .C(n18), .Z(n16) );
  ND2 U103 ( .A(n19), .B(n31), .Z(n17) );
  AO6 U104 ( .A(n19), .B(n32), .C(n20), .Z(n18) );
  AO7 U105 ( .A(n21), .B(n29), .C(n22), .Z(n20) );
  EO U106 ( .A(n23), .B(n2), .Z(SUM[9]) );
  ND2 U107 ( .A(n61), .B(n22), .Z(n2) );
  AO6 U108 ( .A(n24), .B(n44), .C(n25), .Z(n23) );
  IV U109 ( .A(n21), .Z(n61) );
  EO U110 ( .A(n30), .B(n3), .Z(SUM[8]) );
  ND2 U111 ( .A(n62), .B(n29), .Z(n3) );
  AO6 U112 ( .A(n44), .B(n31), .C(n32), .Z(n30) );
  IV U113 ( .A(n26), .Z(n62) );
  AO6 U114 ( .A(n16), .B(n114), .C(n115), .Z(n9) );
  AO7 U115 ( .A(n34), .B(n26), .C(n29), .Z(n25) );
  IV U116 ( .A(n32), .Z(n34) );
  EN U117 ( .A(n44), .B(n5), .Z(SUM[6]) );
  ND2 U118 ( .A(n64), .B(n43), .Z(n5) );
  IV U119 ( .A(n42), .Z(n64) );
  IV U120 ( .A(n43), .Z(n41) );
  AO7 U121 ( .A(n55), .B(n1), .C(n56), .Z(n54) );
  IVP U122 ( .A(n57), .Z(n1) );
  EN U123 ( .A(n8), .B(n57), .Z(SUM[3]) );
  ND2 U124 ( .A(n67), .B(n56), .Z(n8) );
  IV U125 ( .A(n55), .Z(n67) );
  OR2 U126 ( .A(B[0]), .B(A[0]), .Z(n117) );
  EN U127 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  ND2 U128 ( .A(A[8]), .B(B[8]), .Z(n29) );
  ND2 U129 ( .A(A[6]), .B(B[6]), .Z(n43) );
  ND2 U130 ( .A(A[7]), .B(B[7]), .Z(n38) );
  ND2 U131 ( .A(A[3]), .B(B[3]), .Z(n56) );
  ND2 U132 ( .A(A[9]), .B(B[9]), .Z(n22) );
  ND2 U133 ( .A(A[5]), .B(B[5]), .Z(n49) );
  ND2 U134 ( .A(A[4]), .B(B[4]), .Z(n52) );
endmodule


module prime_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] DIFF;
  input CI;
  output CO;
  wire   n3, n4, n9, n10, n11, n13, n14, n15, n16, n17, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n51, n52, n53,
         n55, n58, n59, n60, n61, n62, n64, n65, n68, n70, n71, n72, n76, n77,
         n78, n79, n80, n85, n86, n93, n150, n151, n152, n153, n155, n157,
         n158, n159, n160, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171;
  assign n11 = B[10];
  assign n17 = B[9];
  assign n80 = B[2];
  assign n85 = B[1];
  assign DIFF[0] = n86;
  assign n86 = B[0];

  MUX21LP U4 ( .A(n153), .B(n150), .S(n23), .Z(DIFF[13]) );
  MUX21LP U14 ( .A(n14), .B(n13), .S(n23), .Z(DIFF[12]) );
  NR2 U17 ( .A(n21), .B(n168), .Z(n15) );
  NR2 U18 ( .A(n22), .B(n168), .Z(n16) );
  NR2 U25 ( .A(A[11]), .B(n167), .Z(n21) );
  MUX21LP U28 ( .A(n26), .B(n27), .S(n55), .Z(n23) );
  EOP U50 ( .A(n46), .B(n52), .Z(n43) );
  MUX21LP U51 ( .A(n47), .B(n48), .S(n51), .Z(n44) );
  MUX21LP U52 ( .A(n47), .B(n48), .S(n52), .Z(n45) );
  NR2 U54 ( .A(n169), .B(A[8]), .Z(n47) );
  MUX21LP U64 ( .A(n59), .B(n58), .S(n68), .Z(n55) );
  MUX21LP U67 ( .A(n61), .B(n62), .S(n64), .Z(n58) );
  MUX21LP U68 ( .A(n61), .B(n62), .S(n65), .Z(n59) );
  NR2 U70 ( .A(n164), .B(A[6]), .Z(n61) );
  NR2 U74 ( .A(n93), .B(A[5]), .Z(n64) );
  MUX21LP U79 ( .A(n70), .B(n71), .S(n72), .Z(n68) );
  NR2 U81 ( .A(n170), .B(A[4]), .Z(n70) );
  ENP U117 ( .A(n170), .B(A[4]), .Z(n155) );
  B5I U118 ( .A(n17), .Z(n168) );
  IVA U119 ( .A(n80), .Z(n166) );
  EOP U120 ( .A(n15), .B(n162), .Z(n150) );
  IVP U121 ( .A(n166), .Z(n165) );
  MUX21L U122 ( .A(n4), .B(n3), .S(n23), .Z(DIFF[14]) );
  EOP U123 ( .A(A[11]), .B(n167), .Z(n20) );
  IVAP U124 ( .A(B[3]), .Z(n171) );
  NR2P U125 ( .A(n168), .B(A[9]), .Z(n38) );
  IVP U126 ( .A(B[8]), .Z(n169) );
  IV U127 ( .A(B[7]), .Z(n163) );
  EOP U128 ( .A(n46), .B(n51), .Z(n42) );
  NR2P U129 ( .A(n163), .B(A[7]), .Z(n51) );
  IV U130 ( .A(B[6]), .Z(n164) );
  EOP U131 ( .A(n38), .B(n32), .Z(n28) );
  EOP U132 ( .A(n32), .B(n39), .Z(n29) );
  ENP U133 ( .A(n85), .B(n86), .Z(DIFF[1]) );
  ENP U134 ( .A(n162), .B(A[10]), .Z(n32) );
  EOP U135 ( .A(n16), .B(n162), .Z(n153) );
  IVP U136 ( .A(n11), .Z(n162) );
  MUX21LP U137 ( .A(n33), .B(n34), .S(n39), .Z(n31) );
  MUX21LP U138 ( .A(n33), .B(n34), .S(n38), .Z(n30) );
  NR2P U139 ( .A(n162), .B(A[10]), .Z(n33) );
  IV U140 ( .A(B[11]), .Z(n167) );
  MUX21L U141 ( .A(n36), .B(n35), .S(n53), .Z(DIFF[9]) );
  IV U142 ( .A(n44), .Z(n40) );
  IV U143 ( .A(n45), .Z(n41) );
  ND2P U144 ( .A(n165), .B(n160), .Z(n79) );
  EO U145 ( .A(n72), .B(n155), .Z(DIFF[4]) );
  MUX21LP U146 ( .A(n43), .B(n42), .S(n53), .Z(DIFF[8]) );
  EOP U147 ( .A(n151), .B(n152), .Z(DIFF[7]) );
  EN U148 ( .A(n163), .B(A[7]), .Z(n152) );
  NR2P U149 ( .A(n171), .B(n86), .Z(n77) );
  IVDA U150 ( .A(n55), .Y(n53), .Z(n151) );
  ND2 U151 ( .A(n164), .B(A[6]), .Z(n62) );
  MUX21L U152 ( .A(n31), .B(n30), .S(n44), .Z(n26) );
  MUX21L U153 ( .A(n31), .B(n30), .S(n45), .Z(n27) );
  ND2 U154 ( .A(n170), .B(A[4]), .Z(n71) );
  EO U155 ( .A(n41), .B(n37), .Z(n36) );
  EO U156 ( .A(n40), .B(n37), .Z(n35) );
  EO U157 ( .A(n168), .B(A[9]), .Z(n37) );
  ND2 U158 ( .A(n168), .B(A[9]), .Z(n39) );
  MUX21L U159 ( .A(n24), .B(n25), .S(n55), .Z(DIFF[10]) );
  MUX21L U160 ( .A(n29), .B(n28), .S(n44), .Z(n24) );
  MUX21L U161 ( .A(n29), .B(n28), .S(n45), .Z(n25) );
  MUX21L U162 ( .A(n157), .B(n158), .S(n68), .Z(DIFF[6]) );
  EN U163 ( .A(n60), .B(n65), .Z(n157) );
  EN U164 ( .A(n64), .B(n60), .Z(n158) );
  EN U165 ( .A(n164), .B(A[6]), .Z(n60) );
  EO U166 ( .A(n166), .B(n160), .Z(DIFF[2]) );
  EOP U167 ( .A(n23), .B(n20), .Z(DIFF[11]) );
  EO U168 ( .A(n68), .B(n159), .Z(DIFF[5]) );
  EO U169 ( .A(n93), .B(A[5]), .Z(n159) );
  MUX21H U170 ( .A(n78), .B(n77), .S(n79), .Z(n72) );
  EO U171 ( .A(n169), .B(A[8]), .Z(n46) );
  ND2 U172 ( .A(n93), .B(A[5]), .Z(n65) );
  ND2 U173 ( .A(n163), .B(A[7]), .Z(n52) );
  ND2 U174 ( .A(n169), .B(A[8]), .Z(n48) );
  AN2P U175 ( .A(n86), .B(n85), .Z(n160) );
  EO U176 ( .A(n76), .B(n79), .Z(DIFF[3]) );
  EO U177 ( .A(n171), .B(n86), .Z(n76) );
  EO U178 ( .A(n10), .B(A[14]), .Z(n4) );
  EO U179 ( .A(n9), .B(A[14]), .Z(n3) );
  EO U180 ( .A(n21), .B(n17), .Z(n13) );
  EO U181 ( .A(n22), .B(n17), .Z(n14) );
  ND2 U182 ( .A(A[11]), .B(n167), .Z(n22) );
  ND2 U183 ( .A(n16), .B(n11), .Z(n10) );
  ND2 U184 ( .A(n15), .B(n11), .Z(n9) );
  ND2 U185 ( .A(n162), .B(A[10]), .Z(n34) );
  IV U186 ( .A(B[5]), .Z(n93) );
  ND2 U187 ( .A(n171), .B(n86), .Z(n78) );
  IVA U188 ( .A(B[4]), .Z(n170) );
endmodule


module prime_DW01_add_112 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n36,
         n37, n38, n39, n40, n41, n44, n45, n46, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n68, n69,
         n70, n71, n72, n73, n74, n123, n124, n125, n126, n127;

  NR2 U7 ( .A(n16), .B(n15), .Z(n14) );
  NR2 U10 ( .A(n21), .B(n19), .Z(n17) );
  NR2 U12 ( .A(A[11]), .B(B[11]), .Z(n19) );
  NR2 U14 ( .A(A[10]), .B(B[10]), .Z(n21) );
  NR2 U20 ( .A(n33), .B(n28), .Z(n26) );
  NR2 U28 ( .A(n40), .B(n33), .Z(n31) );
  NR2 U42 ( .A(n49), .B(n44), .Z(n38) );
  NR2 U46 ( .A(A[7]), .B(B[7]), .Z(n44) );
  NR2 U54 ( .A(A[6]), .B(B[6]), .Z(n49) );
  AO6P U58 ( .A(n53), .B(n61), .C(n54), .Z(n52) );
  NR2 U59 ( .A(n58), .B(n55), .Z(n53) );
  NR2 U63 ( .A(A[5]), .B(B[5]), .Z(n55) );
  NR2 U69 ( .A(A[4]), .B(B[4]), .Z(n58) );
  NR2 U77 ( .A(A[3]), .B(B[3]), .Z(n62) );
  FA1A U79 ( .A(n65), .B(A[2]), .CI(B[2]), .CO(n64), .S(SUM[2]) );
  FA1A U80 ( .A(n127), .B(A[1]), .CI(B[1]), .CO(n65), .S(SUM[1]) );
  AN2 U88 ( .A(n18), .B(n14), .Z(n123) );
  AN2 U89 ( .A(n17), .B(n14), .Z(n124) );
  AN2P U90 ( .A(n125), .B(n126), .Z(n28) );
  IV U91 ( .A(A[9]), .Z(n125) );
  IVDA U92 ( .A(B[9]), .Y(n126) );
  AO7P U93 ( .A(n52), .B(n24), .C(n25), .Z(n23) );
  ENP U94 ( .A(n8), .B(n64), .Z(SUM[3]) );
  IV U95 ( .A(n39), .Z(n41) );
  AO6P U96 ( .A(n23), .B(n124), .C(n123), .Z(n9) );
  IV U97 ( .A(n38), .Z(n40) );
  IV U98 ( .A(n50), .Z(n48) );
  AO6P U99 ( .A(n26), .B(n39), .C(n27), .Z(n25) );
  IV U100 ( .A(n61), .Z(n60) );
  AO7 U101 ( .A(n44), .B(n50), .C(n45), .Z(n39) );
  IV U102 ( .A(n9), .Z(CO) );
  AO7 U103 ( .A(n28), .B(n36), .C(n29), .Z(n27) );
  AO7 U104 ( .A(n41), .B(n33), .C(n36), .Z(n32) );
  ND2 U105 ( .A(A[9]), .B(B[9]), .Z(n29) );
  EO U106 ( .A(n30), .B(n2), .Z(SUM[9]) );
  ND2 U107 ( .A(n68), .B(n29), .Z(n2) );
  AO6 U108 ( .A(n31), .B(n51), .C(n32), .Z(n30) );
  IV U109 ( .A(n28), .Z(n68) );
  EO U110 ( .A(n37), .B(n3), .Z(SUM[8]) );
  ND2 U111 ( .A(n69), .B(n36), .Z(n3) );
  AO6 U112 ( .A(n51), .B(n38), .C(n39), .Z(n37) );
  IV U113 ( .A(n33), .Z(n69) );
  EO U114 ( .A(n46), .B(n4), .Z(SUM[7]) );
  ND2 U115 ( .A(n70), .B(n45), .Z(n4) );
  AO6 U116 ( .A(n51), .B(n71), .C(n48), .Z(n46) );
  IV U117 ( .A(n44), .Z(n70) );
  IV U118 ( .A(n49), .Z(n71) );
  ND2 U119 ( .A(n71), .B(n50), .Z(n5) );
  ND2 U120 ( .A(n38), .B(n26), .Z(n24) );
  ND2 U121 ( .A(A[6]), .B(B[6]), .Z(n50) );
  ND2 U122 ( .A(A[8]), .B(B[8]), .Z(n36) );
  ND2 U123 ( .A(A[7]), .B(B[7]), .Z(n45) );
  IV U124 ( .A(n52), .Z(n51) );
  AO7 U125 ( .A(n19), .B(n22), .C(n20), .Z(n18) );
  ND2 U126 ( .A(A[10]), .B(B[10]), .Z(n22) );
  EN U127 ( .A(n57), .B(n6), .Z(SUM[5]) );
  EN U128 ( .A(n51), .B(n5), .Z(SUM[6]) );
  ND2 U129 ( .A(n72), .B(n56), .Z(n6) );
  EO U130 ( .A(n7), .B(n60), .Z(SUM[4]) );
  ND2 U131 ( .A(n73), .B(n59), .Z(n7) );
  IVDA U132 ( .A(B[14]), .Y(n15) );
  ND2 U133 ( .A(B[12]), .B(B[13]), .Z(n16) );
  AO7 U134 ( .A(n62), .B(n1), .C(n63), .Z(n61) );
  IVP U135 ( .A(n64), .Z(n1) );
  ND2 U136 ( .A(n74), .B(n63), .Z(n8) );
  IV U137 ( .A(n62), .Z(n74) );
  OR2 U138 ( .A(B[0]), .B(A[0]), .Z(n127) );
  EN U139 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AO7 U140 ( .A(n60), .B(n58), .C(n59), .Z(n57) );
  IV U141 ( .A(n58), .Z(n73) );
  AO7 U142 ( .A(n55), .B(n59), .C(n56), .Z(n54) );
  IV U143 ( .A(n55), .Z(n72) );
  ND2 U144 ( .A(A[11]), .B(B[11]), .Z(n20) );
  ND2 U145 ( .A(A[5]), .B(B[5]), .Z(n56) );
  NR2P U146 ( .A(A[8]), .B(B[8]), .Z(n33) );
  ND2 U147 ( .A(A[4]), .B(B[4]), .Z(n59) );
  ND2 U148 ( .A(A[3]), .B(B[3]), .Z(n63) );
endmodule


module prime_DW01_add_148 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1, n5, n6, n11, n13, n16, n17, n18, n19, n20, n22, n23, n26, n28,
         n29, n30, n31, n78, n79, n80, n82, n83, n84, n86, n87;

  NR2 U1 ( .A(n13), .B(n78), .Z(CO) );
  NR2 U6 ( .A(n80), .B(n11), .Z(n6) );
  NR2 U20 ( .A(A[5]), .B(B[5]), .Z(n19) );
  MUX21LP U29 ( .A(n28), .B(n29), .S(n1), .Z(n26) );
  NR2 U31 ( .A(A[3]), .B(B[3]), .Z(n28) );
  FA1A U34 ( .A(B[2]), .B(A[2]), .CI(n31), .CO(n30), .S(SUM[2]) );
  FA1AP U43 ( .A(B[1]), .B(A[1]), .CI(n84), .CO(n31), .S(SUM[1]) );
  IVP U44 ( .A(n30), .Z(n1) );
  OR2 U45 ( .A(n5), .B(n87), .Z(n78) );
  ENP U46 ( .A(n22), .B(n18), .Z(n83) );
  NR2P U47 ( .A(A[4]), .B(B[4]), .Z(n22) );
  ENP U48 ( .A(A[5]), .B(B[5]), .Z(n18) );
  EOP U49 ( .A(A[4]), .B(B[4]), .Z(n79) );
  OR2P U50 ( .A(B[0]), .B(A[0]), .Z(n84) );
  MUX21L U51 ( .A(n19), .B(n20), .S(n22), .Z(n16) );
  MUX21L U52 ( .A(n19), .B(n20), .S(n23), .Z(n17) );
  MUX21L U53 ( .A(n17), .B(n16), .S(n26), .Z(n13) );
  EO U54 ( .A(n26), .B(n79), .Z(SUM[4]) );
  ND2 U55 ( .A(B[8]), .B(B[9]), .Z(n80) );
  MUX21L U56 ( .A(n82), .B(n83), .S(n26), .Z(SUM[5]) );
  EN U57 ( .A(n18), .B(n23), .Z(n82) );
  ND2 U58 ( .A(A[3]), .B(B[3]), .Z(n29) );
  EO U59 ( .A(n86), .B(n1), .Z(SUM[3]) );
  EN U60 ( .A(A[3]), .B(B[3]), .Z(n86) );
  EN U61 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  ND2 U62 ( .A(B[6]), .B(B[7]), .Z(n11) );
  ND2 U63 ( .A(n6), .B(B[10]), .Z(n5) );
  ND2 U64 ( .A(A[5]), .B(B[5]), .Z(n20) );
  ND2 U65 ( .A(A[4]), .B(B[4]), .Z(n23) );
  IV U66 ( .A(B[11]), .Z(n87) );
endmodule


module prime_DW01_add_154 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n22, n24, n25, n26, n30, n33, n34, n35, n36, n37, n81,
         n82, n84;

  NR2 U3 ( .A(n3), .B(n4), .Z(n2) );
  AO6P U11 ( .A(n12), .B(n22), .C(n13), .Z(n9) );
  EOP U19 ( .A(n81), .B(n17), .Z(SUM[4]) );
  NR2 U21 ( .A(A[4]), .B(B[4]), .Z(n18) );
  AO7P U26 ( .A(n24), .B(n26), .C(n25), .Z(n22) );
  NR2 U28 ( .A(A[3]), .B(B[3]), .Z(n24) );
  AO7P U39 ( .A(n35), .B(n37), .C(n36), .Z(n33) );
  NR2 U44 ( .A(B[0]), .B(A[0]), .Z(n37) );
  MUX21H U49 ( .A(n11), .B(n10), .S(n82), .Z(SUM[5]) );
  ENP U50 ( .A(B[1]), .B(A[1]), .Z(n34) );
  NR2 U51 ( .A(B[1]), .B(A[1]), .Z(n35) );
  AO5P U52 ( .A(A[2]), .B(B[2]), .C(n33), .Z(n26) );
  NR2P U53 ( .A(n6), .B(n7), .Z(n5) );
  ND2P U54 ( .A(B[9]), .B(B[8]), .Z(n6) );
  IVDA U55 ( .A(n22), .Y(n81), .Z(n82) );
  NR2P U56 ( .A(B[5]), .B(A[5]), .Z(n15) );
  ENP U57 ( .A(B[5]), .B(A[5]), .Z(n14) );
  ND2 U58 ( .A(B[6]), .B(B[7]), .Z(n7) );
  ND2 U59 ( .A(B[11]), .B(B[10]), .Z(n4) );
  IV U60 ( .A(B[12]), .Z(n3) );
  EO U61 ( .A(n14), .B(n19), .Z(n11) );
  EO U62 ( .A(n14), .B(n18), .Z(n10) );
  EN U63 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  EO U64 ( .A(n30), .B(n33), .Z(SUM[2]) );
  ND2 U65 ( .A(A[3]), .B(B[3]), .Z(n25) );
  EN U66 ( .A(A[4]), .B(B[4]), .Z(n17) );
  ND2 U67 ( .A(A[4]), .B(B[4]), .Z(n19) );
  ND2 U68 ( .A(B[1]), .B(A[1]), .Z(n36) );
  EO U69 ( .A(n26), .B(n84), .Z(SUM[3]) );
  EN U70 ( .A(A[3]), .B(B[3]), .Z(n84) );
  EO U71 ( .A(B[2]), .B(A[2]), .Z(n30) );
  EO U72 ( .A(n34), .B(n37), .Z(SUM[1]) );
  AO7 U73 ( .A(n15), .B(n19), .C(n16), .Z(n13) );
  AO7 U74 ( .A(n15), .B(n18), .C(n16), .Z(n12) );
  NR2P U75 ( .A(n1), .B(n9), .Z(CO) );
  ND2 U76 ( .A(n5), .B(n2), .Z(n1) );
  ND2 U77 ( .A(B[5]), .B(A[5]), .Z(n16) );
endmodule


module prime_DW01_add_167 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n8, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n35, n36, n37, n38,
         n39, n40, n83, n84, n85, n86, n87;

  ENP U9 ( .A(n20), .B(n2), .Z(SUM[5]) );
  AO6P U10 ( .A(n16), .B(n24), .C(n17), .Z(n15) );
  NR2 U11 ( .A(n21), .B(n18), .Z(n16) );
  NR2 U15 ( .A(A[5]), .B(B[5]), .Z(n18) );
  EOP U17 ( .A(n23), .B(n3), .Z(SUM[4]) );
  NR2 U21 ( .A(A[4]), .B(B[4]), .Z(n21) );
  NR2 U28 ( .A(A[3]), .B(B[3]), .Z(n25) );
  EOP U30 ( .A(n5), .B(n31), .Z(SUM[2]) );
  AO7P U32 ( .A(n31), .B(n29), .C(n30), .Z(n28) );
  NR2 U35 ( .A(B[2]), .B(A[2]), .Z(n29) );
  EOP U37 ( .A(n6), .B(n36), .Z(SUM[1]) );
  AO6P U38 ( .A(n87), .B(n1), .C(n33), .Z(n31) );
  ND2P U45 ( .A(B[1]), .B(A[1]), .Z(n35) );
  NR2 U47 ( .A(B[0]), .B(A[0]), .Z(n36) );
  AN2P U52 ( .A(B[13]), .B(B[12]), .Z(n83) );
  AO7 U53 ( .A(n25), .B(n27), .C(n26), .Z(n24) );
  AN2P U54 ( .A(B[10]), .B(B[11]), .Z(n84) );
  AN2P U55 ( .A(B[8]), .B(B[9]), .Z(n85) );
  AN2P U56 ( .A(B[6]), .B(B[7]), .Z(n86) );
  ND4P U57 ( .A(n84), .B(n83), .C(n86), .D(n85), .Z(n8) );
  NR2P U58 ( .A(n8), .B(n15), .Z(CO) );
  IVP U59 ( .A(n28), .Z(n27) );
  EO U60 ( .A(n4), .B(n27), .Z(SUM[3]) );
  ND2 U61 ( .A(n38), .B(n22), .Z(n3) );
  IV U62 ( .A(n35), .Z(n33) );
  IVA U63 ( .A(n36), .Z(n1) );
  IV U64 ( .A(n24), .Z(n23) );
  ND2 U65 ( .A(n87), .B(n35), .Z(n6) );
  AO7 U66 ( .A(n18), .B(n22), .C(n19), .Z(n17) );
  EN U67 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  OR2 U68 ( .A(B[1]), .B(A[1]), .Z(n87) );
  AO7 U69 ( .A(n23), .B(n21), .C(n22), .Z(n20) );
  ND2 U70 ( .A(n37), .B(n19), .Z(n2) );
  IV U71 ( .A(n18), .Z(n37) );
  IV U72 ( .A(n21), .Z(n38) );
  ND2 U73 ( .A(n39), .B(n26), .Z(n4) );
  IV U74 ( .A(n25), .Z(n39) );
  ND2 U75 ( .A(n40), .B(n30), .Z(n5) );
  IV U76 ( .A(n29), .Z(n40) );
  ND2 U77 ( .A(A[4]), .B(B[4]), .Z(n22) );
  ND2 U78 ( .A(A[3]), .B(B[3]), .Z(n26) );
  ND2 U79 ( .A(B[2]), .B(A[2]), .Z(n30) );
  ND2 U80 ( .A(A[5]), .B(B[5]), .Z(n19) );
endmodule


module prime_DW01_add_157 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n33, \A[0] , n74;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  ND2P U4 ( .A(B[13]), .B(B[12]), .Z(n8) );
  NR2 U6 ( .A(n12), .B(n11), .Z(n10) );
  ENP U9 ( .A(n18), .B(n1), .Z(SUM[5]) );
  AO6P U10 ( .A(n14), .B(n22), .C(n15), .Z(n13) );
  NR2 U11 ( .A(n19), .B(n16), .Z(n14) );
  NR2 U21 ( .A(A[4]), .B(B[4]), .Z(n19) );
  NR2 U35 ( .A(B[2]), .B(A[2]), .Z(n27) );
  NR2 U38 ( .A(B[1]), .B(A[1]), .Z(n29) );
  ND2 U43 ( .A(n31), .B(n20), .Z(n2) );
  AO7 U44 ( .A(n27), .B(n29), .C(n28), .Z(n26) );
  ND2 U45 ( .A(n33), .B(n28), .Z(n4) );
  OR2 U46 ( .A(A[3]), .B(B[3]), .Z(n74) );
  ND2P U47 ( .A(A[3]), .B(B[3]), .Z(n24) );
  NR2P U48 ( .A(A[5]), .B(B[5]), .Z(n16) );
  ND2P U49 ( .A(B[10]), .B(B[11]), .Z(n9) );
  AO7P U50 ( .A(n23), .B(n25), .C(n24), .Z(n22) );
  NR2P U51 ( .A(A[3]), .B(B[3]), .Z(n23) );
  IV U52 ( .A(n22), .Z(n21) );
  AO7 U53 ( .A(n16), .B(n20), .C(n17), .Z(n15) );
  AO7 U54 ( .A(n21), .B(n19), .C(n20), .Z(n18) );
  ND2 U55 ( .A(n30), .B(n17), .Z(n1) );
  IV U56 ( .A(n16), .Z(n30) );
  EO U57 ( .A(n4), .B(n29), .Z(SUM[2]) );
  IV U58 ( .A(n27), .Z(n33) );
  ND2 U59 ( .A(B[8]), .B(B[9]), .Z(n11) );
  EO U60 ( .A(n21), .B(n2), .Z(SUM[4]) );
  IV U61 ( .A(n19), .Z(n31) );
  EO U62 ( .A(n3), .B(n25), .Z(SUM[3]) );
  ND2 U63 ( .A(n74), .B(n24), .Z(n3) );
  EN U64 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  ND2 U65 ( .A(B[6]), .B(B[7]), .Z(n12) );
  ND2 U66 ( .A(A[4]), .B(B[4]), .Z(n20) );
  ND2 U67 ( .A(B[2]), .B(A[2]), .Z(n28) );
  NR2P U68 ( .A(n9), .B(n8), .Z(n7) );
  NR2P U69 ( .A(n6), .B(n13), .Z(CO) );
  ND2 U70 ( .A(n7), .B(n10), .Z(n6) );
  ND2 U71 ( .A(A[5]), .B(B[5]), .Z(n17) );
  IVAP U72 ( .A(n26), .Z(n25) );
endmodule


module prime_DW01_add_156 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n9, n14, n15, n16, n17, n20, n21, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n41, n42,
         n45, n47, n48, n49, \A[0] , \A[1] , n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n104, n105, n106;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];

  MUX21LP U1 ( .A(n1), .B(n2), .S(n32), .Z(CO) );
  NR2 U17 ( .A(A[8]), .B(B[8]), .Z(n15) );
  MUX21LP U28 ( .A(n27), .B(n28), .S(n31), .Z(n25) );
  MUX21LP U37 ( .A(n36), .B(n35), .S(n45), .Z(n32) );
  MUX21LP U52 ( .A(n47), .B(n48), .S(n49), .Z(n45) );
  NR2 U57 ( .A(B[2]), .B(A[2]), .Z(n49) );
  ENP U62 ( .A(n17), .B(n14), .Z(SUM[8]) );
  EO U63 ( .A(n37), .B(n42), .Z(n34) );
  MUX21L U64 ( .A(n38), .B(n39), .S(n42), .Z(n36) );
  IVDA U65 ( .A(A[4]), .Z(n94) );
  NR2P U66 ( .A(A[3]), .B(B[3]), .Z(n47) );
  NR2 U67 ( .A(n94), .B(B[4]), .Z(n95) );
  NR2P U68 ( .A(n16), .B(n105), .Z(n4) );
  ND2P U69 ( .A(A[4]), .B(B[4]), .Z(n42) );
  IVDA U70 ( .A(A[6]), .Z(n96) );
  B2I U71 ( .A(n32), .Z2(n97) );
  NR2P U72 ( .A(A[7]), .B(B[7]), .Z(n27) );
  EOP U73 ( .A(n94), .B(B[4]), .Z(n102) );
  ND2 U74 ( .A(A[5]), .B(B[5]), .Z(n39) );
  NR2 U75 ( .A(A[5]), .B(B[5]), .Z(n98) );
  NR2P U76 ( .A(n15), .B(n105), .Z(n3) );
  EOP U77 ( .A(A[5]), .B(B[5]), .Z(n37) );
  NR2 U78 ( .A(A[5]), .B(B[5]), .Z(n38) );
  NR2P U79 ( .A(A[6]), .B(B[6]), .Z(n30) );
  ND2P U80 ( .A(A[6]), .B(B[6]), .Z(n31) );
  NR2 U81 ( .A(n96), .B(B[6]), .Z(n99) );
  ENP U82 ( .A(n26), .B(n99), .Z(n101) );
  MUX21L U83 ( .A(n27), .B(n28), .S(n30), .Z(n24) );
  IV U84 ( .A(n25), .Z(n21) );
  IV U85 ( .A(n24), .Z(n20) );
  EN U86 ( .A(n26), .B(n31), .Z(n100) );
  EN U87 ( .A(A[7]), .B(B[7]), .Z(n26) );
  EO U88 ( .A(n45), .B(n102), .Z(SUM[4]) );
  EOP U89 ( .A(n104), .B(n49), .Z(SUM[3]) );
  EN U90 ( .A(A[3]), .B(B[3]), .Z(n104) );
  ND2 U91 ( .A(A[3]), .B(B[3]), .Z(n48) );
  ND2 U92 ( .A(A[8]), .B(B[8]), .Z(n16) );
  MUX21L U93 ( .A(n101), .B(n100), .S(n97), .Z(SUM[7]) );
  EN U94 ( .A(A[8]), .B(B[8]), .Z(n14) );
  EO U95 ( .A(n97), .B(n29), .Z(SUM[6]) );
  EN U96 ( .A(n96), .B(B[6]), .Z(n29) );
  AN2P U97 ( .A(B[9]), .B(B[10]), .Z(n9) );
  ND2 U98 ( .A(n106), .B(B[12]), .Z(n105) );
  AN2P U99 ( .A(n9), .B(B[11]), .Z(n106) );
  EN U100 ( .A(B[2]), .B(A[2]), .Z(SUM[2]) );
  MUX21L U101 ( .A(n34), .B(n33), .S(n45), .Z(SUM[5]) );
  EO U102 ( .A(n37), .B(n95), .Z(n33) );
  MUX21L U103 ( .A(n20), .B(n21), .S(n97), .Z(n17) );
  MUX21L U104 ( .A(n4), .B(n3), .S(n25), .Z(n2) );
  MUX21L U105 ( .A(n4), .B(n3), .S(n24), .Z(n1) );
  MUX21L U106 ( .A(n98), .B(n39), .S(n41), .Z(n35) );
  ND2 U107 ( .A(A[7]), .B(B[7]), .Z(n28) );
  NR2P U108 ( .A(A[4]), .B(B[4]), .Z(n41) );
endmodule


module prime_DW01_add_176 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n6, n8, n10, n11, n12, n13, n14, n15, n16, n18, n20, n21,
         n23, n25, n26, n27, n29, n31, n32, n33, n81, n82, n83, n84, n85, n86,
         n87;

  ND2P U4 ( .A(B[12]), .B(B[13]), .Z(n8) );
  NR2 U7 ( .A(n13), .B(n12), .Z(n11) );
  EOP U10 ( .A(n21), .B(n2), .Z(SUM[5]) );
  MUX21LP U30 ( .A(n29), .B(n84), .S(n32), .Z(n27) );
  FA1A U37 ( .A(n33), .B(A[2]), .CI(B[2]), .CO(n32), .S(SUM[2]) );
  FA1A U38 ( .A(n83), .B(A[1]), .CI(B[1]), .CO(n33), .S(SUM[1]) );
  ENP U46 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  IVA U47 ( .A(n27), .Z(n26) );
  IVA U48 ( .A(n25), .Z(n23) );
  OR2P U49 ( .A(A[5]), .B(B[5]), .Z(n81) );
  IVP U50 ( .A(n20), .Z(n18) );
  ND2 U51 ( .A(n81), .B(n20), .Z(n2) );
  OR2P U52 ( .A(A[4]), .B(B[4]), .Z(n82) );
  IV U53 ( .A(n31), .Z(n29) );
  EN U54 ( .A(n4), .B(n32), .Z(SUM[3]) );
  MUX21L U55 ( .A(n23), .B(n82), .S(n26), .Z(n21) );
  ND2 U56 ( .A(n11), .B(n14), .Z(n10) );
  MUX21L U57 ( .A(n15), .B(n16), .S(n27), .Z(n14) );
  MUX21L U58 ( .A(n18), .B(n81), .S(n82), .Z(n15) );
  MUX21L U59 ( .A(n18), .B(n81), .S(n23), .Z(n16) );
  ND2 U60 ( .A(B[7]), .B(B[6]), .Z(n13) );
  ND2 U61 ( .A(B[8]), .B(B[9]), .Z(n12) );
  ND2 U62 ( .A(n82), .B(n25), .Z(n3) );
  EN U63 ( .A(n3), .B(n26), .Z(SUM[4]) );
  OR2 U64 ( .A(B[0]), .B(A[0]), .Z(n83) );
  ND2 U65 ( .A(n84), .B(n31), .Z(n4) );
  OR2 U66 ( .A(A[3]), .B(B[3]), .Z(n84) );
  ND2 U67 ( .A(A[3]), .B(B[3]), .Z(n31) );
  IV U68 ( .A(B[14]), .Z(n85) );
  ND2P U69 ( .A(n86), .B(n87), .Z(n6) );
  AN2 U70 ( .A(B[11]), .B(B[10]), .Z(n86) );
  NR2P U71 ( .A(n8), .B(n85), .Z(n87) );
  NR2P U72 ( .A(n6), .B(n10), .Z(CO) );
  ND2 U73 ( .A(A[5]), .B(B[5]), .Z(n20) );
  ND2 U74 ( .A(A[4]), .B(B[4]), .Z(n25) );
endmodule


module prime_DW01_add_198 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n7, n10, n12, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n28, n30, n31, n32, n33, n34, n35, n36,
         n37, n39, n81, n82, n83, n84, n85;

  ENP U9 ( .A(n19), .B(n1), .Z(SUM[5]) );
  NR2 U11 ( .A(n17), .B(n20), .Z(n15) );
  EOP U17 ( .A(n22), .B(n2), .Z(SUM[4]) );
  NR2 U21 ( .A(A[4]), .B(B[4]), .Z(n20) );
  AO7P U25 ( .A(n26), .B(n24), .C(n25), .Z(n23) );
  NR2 U28 ( .A(A[3]), .B(B[3]), .Z(n24) );
  AO6P U31 ( .A(n85), .B(n31), .C(n28), .Z(n26) );
  NR2 U42 ( .A(B[1]), .B(A[1]), .Z(n32) );
  NR2 U45 ( .A(B[0]), .B(A[0]), .Z(n34) );
  ND2 U50 ( .A(n36), .B(n21), .Z(n2) );
  ND2 U51 ( .A(n37), .B(n25), .Z(n3) );
  ND2 U52 ( .A(n39), .B(n33), .Z(n5) );
  AN2P U53 ( .A(B[13]), .B(B[12]), .Z(n81) );
  AN2P U54 ( .A(B[6]), .B(B[7]), .Z(n82) );
  ND2 U55 ( .A(B[11]), .B(B[10]), .Z(n10) );
  AO7P U56 ( .A(n17), .B(n21), .C(n18), .Z(n16) );
  ND4P U57 ( .A(n83), .B(n82), .C(n81), .D(n84), .Z(n7) );
  IVA U58 ( .A(n12), .Z(n83) );
  IVA U59 ( .A(n10), .Z(n84) );
  AO6P U60 ( .A(n15), .B(n23), .C(n16), .Z(n14) );
  ND2P U61 ( .A(B[2]), .B(A[2]), .Z(n30) );
  NR2P U62 ( .A(B[5]), .B(A[5]), .Z(n17) );
  EN U63 ( .A(n4), .B(n31), .Z(SUM[2]) );
  AO7 U64 ( .A(n32), .B(n34), .C(n33), .Z(n31) );
  ND2 U65 ( .A(n35), .B(n18), .Z(n1) );
  IV U66 ( .A(n23), .Z(n22) );
  EO U67 ( .A(n5), .B(n34), .Z(SUM[1]) );
  IV U68 ( .A(n32), .Z(n39) );
  IVP U69 ( .A(n30), .Z(n28) );
  IV U70 ( .A(n20), .Z(n36) );
  AO7 U71 ( .A(n22), .B(n20), .C(n21), .Z(n19) );
  EN U72 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  ND2 U73 ( .A(B[1]), .B(A[1]), .Z(n33) );
  EO U74 ( .A(n3), .B(n26), .Z(SUM[3]) );
  IV U75 ( .A(n24), .Z(n37) );
  ND2 U76 ( .A(n85), .B(n30), .Z(n4) );
  OR2 U77 ( .A(B[2]), .B(A[2]), .Z(n85) );
  ND2 U78 ( .A(A[4]), .B(B[4]), .Z(n21) );
  ND2 U79 ( .A(A[3]), .B(B[3]), .Z(n25) );
  IV U80 ( .A(n17), .Z(n35) );
  ND2 U81 ( .A(B[9]), .B(B[8]), .Z(n12) );
  NR2P U82 ( .A(n7), .B(n14), .Z(CO) );
  ND2 U83 ( .A(B[5]), .B(A[5]), .Z(n18) );
endmodule


module prime_DW01_add_204 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n12, n13, n14, n15, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n39, n40, n43, n45, n46, n47, n48, n99, n101, n102, n103, n104;

  NR2 U4 ( .A(n13), .B(n102), .Z(n4) );
  NR2 U5 ( .A(n14), .B(n102), .Z(n5) );
  NR2 U14 ( .A(A[8]), .B(B[8]), .Z(n13) );
  NR2 U27 ( .A(A[7]), .B(B[7]), .Z(n25) );
  NR2 U31 ( .A(A[6]), .B(B[6]), .Z(n28) );
  MUX21LP U34 ( .A(n34), .B(n33), .S(n43), .Z(n30) );
  NR2 U40 ( .A(A[5]), .B(B[5]), .Z(n36) );
  NR2 U44 ( .A(A[4]), .B(B[4]), .Z(n39) );
  NR2 U51 ( .A(A[3]), .B(B[3]), .Z(n45) );
  FA1A U55 ( .A(B[1]), .B(A[1]), .CI(n104), .CO(n48), .S(SUM[1]) );
  ENP U63 ( .A(A[3]), .B(B[3]), .Z(n101) );
  IVP U64 ( .A(n47), .Z(n1) );
  EOP U65 ( .A(A[5]), .B(B[5]), .Z(n35) );
  ENP U66 ( .A(A[6]), .B(B[6]), .Z(n27) );
  FA1AP U67 ( .A(B[2]), .B(A[2]), .CI(n48), .CO(n47), .S(SUM[2]) );
  MUX21LP U68 ( .A(n25), .B(n26), .S(n29), .Z(n23) );
  EO U69 ( .A(n30), .B(n27), .Z(SUM[6]) );
  MUX21L U70 ( .A(n18), .B(n19), .S(n30), .Z(n15) );
  MUX21L U71 ( .A(n2), .B(n3), .S(n30), .Z(CO) );
  ENP U72 ( .A(A[8]), .B(B[8]), .Z(n12) );
  ENP U73 ( .A(A[7]), .B(B[7]), .Z(n24) );
  EOP U74 ( .A(A[4]), .B(B[4]), .Z(n99) );
  IV U75 ( .A(n23), .Z(n19) );
  MUX21LP U76 ( .A(n25), .B(n26), .S(n28), .Z(n22) );
  ENP U77 ( .A(n15), .B(n12), .Z(SUM[8]) );
  OR2P U78 ( .A(B[0]), .B(A[0]), .Z(n104) );
  IVP U79 ( .A(n22), .Z(n18) );
  EO U80 ( .A(n24), .B(n29), .Z(n21) );
  MUX21H U81 ( .A(n20), .B(n21), .S(n30), .Z(SUM[7]) );
  EO U82 ( .A(n28), .B(n24), .Z(n20) );
  MUX21L U83 ( .A(n36), .B(n37), .S(n40), .Z(n34) );
  MUX21L U84 ( .A(n36), .B(n37), .S(n39), .Z(n33) );
  MUX21L U85 ( .A(n45), .B(n46), .S(n1), .Z(n43) );
  MUX21L U86 ( .A(n5), .B(n4), .S(n23), .Z(n3) );
  MUX21L U87 ( .A(n5), .B(n4), .S(n22), .Z(n2) );
  ND2 U88 ( .A(A[8]), .B(B[8]), .Z(n14) );
  MUX21L U89 ( .A(n32), .B(n31), .S(n43), .Z(SUM[5]) );
  EO U90 ( .A(n35), .B(n40), .Z(n32) );
  EO U91 ( .A(n39), .B(n35), .Z(n31) );
  EO U92 ( .A(n43), .B(n99), .Z(SUM[4]) );
  EO U93 ( .A(n101), .B(n1), .Z(SUM[3]) );
  ND2 U94 ( .A(n103), .B(B[11]), .Z(n102) );
  AN2P U95 ( .A(B[10]), .B(B[9]), .Z(n103) );
  EN U96 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  ND2 U97 ( .A(A[6]), .B(B[6]), .Z(n29) );
  ND2 U98 ( .A(A[3]), .B(B[3]), .Z(n46) );
  ND2 U99 ( .A(A[5]), .B(B[5]), .Z(n37) );
  ND2 U100 ( .A(A[4]), .B(B[4]), .Z(n40) );
  ND2 U101 ( .A(A[7]), .B(B[7]), .Z(n26) );
endmodule


module prime_DW01_add_201 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n12, n13, n14, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n42, n43, n44, n45, n46, n47, n95, n97, n98;

  NR2 U4 ( .A(n12), .B(n97), .Z(n4) );
  NR2 U5 ( .A(n13), .B(n97), .Z(n5) );
  ENP U10 ( .A(n14), .B(n95), .Z(SUM[8]) );
  NR2 U13 ( .A(A[8]), .B(B[8]), .Z(n12) );
  NR2 U26 ( .A(A[7]), .B(B[7]), .Z(n24) );
  EOP U34 ( .A(n38), .B(n34), .Z(n30) );
  NR2 U39 ( .A(A[5]), .B(B[5]), .Z(n35) );
  MUX21LP U48 ( .A(n44), .B(n45), .S(n1), .Z(n42) );
  NR2 U50 ( .A(A[3]), .B(B[3]), .Z(n44) );
  FA1 U62 ( .A(B[1]), .B(A[1]), .CI(n98), .CO(n47), .S(SUM[1]) );
  ENP U63 ( .A(A[4]), .B(B[4]), .Z(n37) );
  MUX21L U64 ( .A(n35), .B(n36), .S(n39), .Z(n33) );
  EN U65 ( .A(n42), .B(n37), .Z(SUM[4]) );
  NR2P U66 ( .A(A[4]), .B(B[4]), .Z(n38) );
  EOP U67 ( .A(A[3]), .B(B[3]), .Z(n43) );
  NR2P U68 ( .A(A[6]), .B(B[6]), .Z(n27) );
  EOP U69 ( .A(n27), .B(n23), .Z(n19) );
  MUX21L U70 ( .A(n24), .B(n25), .S(n27), .Z(n21) );
  EOP U71 ( .A(n34), .B(n39), .Z(n31) );
  ENP U72 ( .A(A[6]), .B(B[6]), .Z(n26) );
  EOP U73 ( .A(A[5]), .B(B[5]), .Z(n34) );
  MUX21LP U74 ( .A(n33), .B(n32), .S(n42), .Z(n29) );
  IV U75 ( .A(n21), .Z(n17) );
  MUX21LP U76 ( .A(n24), .B(n25), .S(n28), .Z(n22) );
  MUX21LP U77 ( .A(n2), .B(n3), .S(n29), .Z(CO) );
  EN U78 ( .A(A[8]), .B(B[8]), .Z(n95) );
  OR2P U79 ( .A(B[0]), .B(A[0]), .Z(n98) );
  MUX21L U80 ( .A(n31), .B(n30), .S(n42), .Z(SUM[5]) );
  MUX21L U81 ( .A(n35), .B(n36), .S(n38), .Z(n32) );
  ND2 U82 ( .A(A[4]), .B(B[4]), .Z(n39) );
  IVP U83 ( .A(n22), .Z(n18) );
  EN U84 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  MUX21L U85 ( .A(n5), .B(n4), .S(n22), .Z(n3) );
  MUX21L U86 ( .A(n5), .B(n4), .S(n21), .Z(n2) );
  MUX21H U87 ( .A(n19), .B(n20), .S(n29), .Z(SUM[7]) );
  EO U88 ( .A(n23), .B(n28), .Z(n20) );
  EN U89 ( .A(A[7]), .B(B[7]), .Z(n23) );
  EO U90 ( .A(n29), .B(n26), .Z(SUM[6]) );
  ENP U91 ( .A(n43), .B(n1), .Z(SUM[3]) );
  MUX21L U92 ( .A(n17), .B(n18), .S(n29), .Z(n14) );
  ND2 U93 ( .A(A[8]), .B(B[8]), .Z(n13) );
  ND2 U94 ( .A(B[9]), .B(B[10]), .Z(n97) );
  ND2 U95 ( .A(A[5]), .B(B[5]), .Z(n36) );
  FA1A U96 ( .A(B[2]), .B(A[2]), .CI(n47), .CO(n46), .S(SUM[2]) );
  IVP U97 ( .A(n46), .Z(n1) );
  ND2 U98 ( .A(A[3]), .B(B[3]), .Z(n45) );
  ND2 U99 ( .A(A[7]), .B(B[7]), .Z(n25) );
  ND2 U100 ( .A(A[6]), .B(B[6]), .Z(n28) );
endmodule


module prime_DW01_add_205 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n11, n17, n18, n19, n22, n23, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n47, n49, n50, n51, n52, n100, n101, n102, n103, n104, n106,
         n107;

  NR2 U4 ( .A(n17), .B(n103), .Z(n5) );
  NR2 U5 ( .A(n18), .B(n103), .Z(n6) );
  NR2 U17 ( .A(A[8]), .B(B[8]), .Z(n17) );
  EOP U32 ( .A(n34), .B(n31), .Z(SUM[6]) );
  MUX21LP U37 ( .A(n38), .B(n37), .S(n47), .Z(n34) );
  MUX21LP U52 ( .A(n49), .B(n50), .S(n1), .Z(n47) );
  NR2 U54 ( .A(A[3]), .B(B[3]), .Z(n49) );
  FA1A U57 ( .A(B[2]), .B(A[2]), .CI(n52), .CO(n51), .S(SUM[2]) );
  FA1A U58 ( .A(n107), .B(A[1]), .CI(B[1]), .CO(n52), .S(SUM[1]) );
  MUX21L U66 ( .A(n29), .B(n30), .S(n32), .Z(n26) );
  EOP U67 ( .A(n19), .B(n101), .Z(SUM[8]) );
  ENP U68 ( .A(n28), .B(n33), .Z(n100) );
  ND2P U69 ( .A(A[4]), .B(B[4]), .Z(n44) );
  ENP U70 ( .A(A[4]), .B(B[4]), .Z(n42) );
  EN U71 ( .A(n47), .B(n42), .Z(SUM[4]) );
  MUX21L U72 ( .A(n40), .B(n41), .S(n43), .Z(n37) );
  MUX21L U73 ( .A(n40), .B(n41), .S(n44), .Z(n38) );
  NR2P U74 ( .A(A[5]), .B(B[5]), .Z(n40) );
  AN2P U75 ( .A(B[9]), .B(B[10]), .Z(n11) );
  MUX21L U76 ( .A(n29), .B(n30), .S(n33), .Z(n27) );
  ND2P U77 ( .A(A[6]), .B(B[6]), .Z(n33) );
  NR2P U78 ( .A(A[7]), .B(B[7]), .Z(n29) );
  EOP U79 ( .A(n39), .B(n44), .Z(n36) );
  ENP U80 ( .A(A[6]), .B(B[6]), .Z(n31) );
  NR2P U81 ( .A(A[4]), .B(B[4]), .Z(n43) );
  EOP U82 ( .A(n43), .B(n39), .Z(n35) );
  NR2P U83 ( .A(A[6]), .B(B[6]), .Z(n32) );
  EOP U84 ( .A(A[5]), .B(B[5]), .Z(n39) );
  IV U85 ( .A(n26), .Z(n22) );
  MUX21LP U86 ( .A(n3), .B(n4), .S(n34), .Z(CO) );
  EO U87 ( .A(A[8]), .B(B[8]), .Z(n101) );
  IVP U88 ( .A(n27), .Z(n23) );
  MUX21L U89 ( .A(n22), .B(n23), .S(n34), .Z(n19) );
  MUX21L U90 ( .A(n6), .B(n5), .S(n27), .Z(n4) );
  MUX21L U91 ( .A(n6), .B(n5), .S(n26), .Z(n3) );
  MUX21L U92 ( .A(n102), .B(n100), .S(n34), .Z(SUM[7]) );
  ND2 U93 ( .A(A[8]), .B(B[8]), .Z(n18) );
  EN U94 ( .A(n32), .B(n28), .Z(n102) );
  ND2 U95 ( .A(n104), .B(B[12]), .Z(n103) );
  AN2P U96 ( .A(n11), .B(B[11]), .Z(n104) );
  MUX21L U97 ( .A(n36), .B(n35), .S(n47), .Z(SUM[5]) );
  EN U98 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  EN U99 ( .A(A[7]), .B(B[7]), .Z(n28) );
  ND2 U100 ( .A(A[3]), .B(B[3]), .Z(n50) );
  EOP U101 ( .A(n106), .B(n1), .Z(SUM[3]) );
  EN U102 ( .A(A[3]), .B(B[3]), .Z(n106) );
  IVP U103 ( .A(n51), .Z(n1) );
  OR2 U104 ( .A(B[0]), .B(A[0]), .Z(n107) );
  ND2 U105 ( .A(A[5]), .B(B[5]), .Z(n41) );
  ND2 U106 ( .A(A[7]), .B(B[7]), .Z(n30) );
endmodule


module prime_DW01_add_203 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n12, n13, n14, n15, n18, n19, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n43, n44, n45, n46, n47, \A[0] , n95, n96, n97, n98, n100, n101,
         n102, n103, n104;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  MUX21LP U1 ( .A(n2), .B(n3), .S(n30), .Z(CO) );
  NR2 U4 ( .A(n13), .B(n102), .Z(n4) );
  NR2 U5 ( .A(n14), .B(n102), .Z(n5) );
  NR2 U14 ( .A(A[8]), .B(B[8]), .Z(n13) );
  MUX21LP U34 ( .A(n34), .B(n33), .S(n43), .Z(n30) );
  ND2P U45 ( .A(A[4]), .B(B[4]), .Z(n40) );
  MUX21LP U49 ( .A(n45), .B(n46), .S(n1), .Z(n43) );
  NR2 U51 ( .A(A[3]), .B(B[3]), .Z(n45) );
  IVDA U62 ( .A(A[4]), .Z(n97) );
  IVP U63 ( .A(n47), .Z(n1) );
  ENP U64 ( .A(n44), .B(n1), .Z(SUM[3]) );
  FA1P U65 ( .A(B[2]), .B(A[2]), .CI(n104), .CO(n47), .S(SUM[2]) );
  B2I U66 ( .A(n33), .Z2(n95) );
  MUX21L U67 ( .A(n36), .B(n37), .S(n39), .Z(n33) );
  MUX21LP U68 ( .A(n34), .B(n95), .S(n43), .Z(n96) );
  EN U69 ( .A(n97), .B(B[4]), .Z(n38) );
  NR2P U70 ( .A(A[7]), .B(B[7]), .Z(n25) );
  NR2 U71 ( .A(n97), .B(B[4]), .Z(n98) );
  EOP U72 ( .A(n96), .B(n27), .Z(SUM[6]) );
  MUX21L U73 ( .A(n18), .B(n19), .S(n96), .Z(n15) );
  MUX21L U74 ( .A(n25), .B(n26), .S(n28), .Z(n22) );
  EOP U75 ( .A(n35), .B(n40), .Z(n32) );
  EOP U76 ( .A(n98), .B(n35), .Z(n31) );
  ENP U77 ( .A(A[6]), .B(B[6]), .Z(n27) );
  ENP U78 ( .A(n29), .B(n24), .Z(n101) );
  MUX21L U79 ( .A(n25), .B(n26), .S(n29), .Z(n23) );
  ENP U80 ( .A(n28), .B(n24), .Z(n100) );
  NR2P U81 ( .A(A[6]), .B(B[6]), .Z(n28) );
  EOP U82 ( .A(A[5]), .B(B[5]), .Z(n35) );
  MUX21L U83 ( .A(n36), .B(n37), .S(n40), .Z(n34) );
  NR2P U84 ( .A(A[5]), .B(B[5]), .Z(n36) );
  IV U85 ( .A(n23), .Z(n19) );
  IV U86 ( .A(n22), .Z(n18) );
  ENP U87 ( .A(n15), .B(n12), .Z(SUM[8]) );
  OR2P U88 ( .A(B[1]), .B(A[1]), .Z(n104) );
  MUX21L U89 ( .A(n32), .B(n31), .S(n43), .Z(SUM[5]) );
  EN U90 ( .A(n43), .B(n38), .Z(SUM[4]) );
  MUX21L U91 ( .A(n100), .B(n101), .S(n96), .Z(SUM[7]) );
  MUX21L U92 ( .A(n5), .B(n4), .S(n23), .Z(n3) );
  MUX21L U93 ( .A(n5), .B(n4), .S(n22), .Z(n2) );
  ND2 U94 ( .A(A[3]), .B(B[3]), .Z(n46) );
  ND2 U95 ( .A(A[8]), .B(B[8]), .Z(n14) );
  EN U96 ( .A(A[8]), .B(B[8]), .Z(n12) );
  EO U97 ( .A(A[3]), .B(B[3]), .Z(n44) );
  EN U98 ( .A(A[7]), .B(B[7]), .Z(n24) );
  ND2 U99 ( .A(n103), .B(B[11]), .Z(n102) );
  AN2P U100 ( .A(B[9]), .B(B[10]), .Z(n103) );
  ND2 U101 ( .A(A[5]), .B(B[5]), .Z(n37) );
  EN U102 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  NR2P U103 ( .A(A[4]), .B(B[4]), .Z(n39) );
  ND2 U104 ( .A(A[7]), .B(B[7]), .Z(n26) );
  ND2 U105 ( .A(A[6]), .B(B[6]), .Z(n29) );
endmodule


module prime_DW01_add_232 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n6, n8, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n40, n41, n50, n51, n54, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n71, n72, n79, n80, n81, n83, n84, n86, n88, n89, n90, \B[0] , \B[1] ,
         n140, n141, n142, n143, n144, n146, n147, n148, n149, n150, n151,
         n152, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166;
  assign n6 = B[11];
  assign n8 = B[10];
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];
  assign SUM[1] = \B[1] ;
  assign \B[1]  = B[1];

  OR2 U1 ( .A(n10), .B(n166), .Z(SUM[14]) );
  MUX21LP U3 ( .A(n155), .B(n142), .S(n10), .Z(SUM[13]) );
  ENP U10 ( .A(n10), .B(A[12]), .Z(SUM[12]) );
  MUX21LP U14 ( .A(n13), .B(n14), .S(n56), .Z(n10) );
  MUX21LP U21 ( .A(n20), .B(n21), .S(n25), .Z(n17) );
  MUX21LP U22 ( .A(n20), .B(n21), .S(n26), .Z(n18) );
  MUX21LP U32 ( .A(n30), .B(n29), .S(n54), .Z(SUM[9]) );
  MUX21LP U38 ( .A(n141), .B(n35), .S(n41), .Z(n32) );
  NR2 U40 ( .A(B[9]), .B(A[9]), .Z(n34) );
  MUX21LP U42 ( .A(n159), .B(n147), .S(n54), .Z(SUM[8]) );
  MUX21LP U48 ( .A(n157), .B(n156), .S(n50), .Z(n41) );
  ENP U82 ( .A(n162), .B(n80), .Z(n72) );
  EOP U89 ( .A(n84), .B(n81), .Z(SUM[4]) );
  MUX21LP U98 ( .A(n88), .B(n89), .S(n90), .Z(n86) );
  NR2 U100 ( .A(B[3]), .B(A[3]), .Z(n88) );
  ENP U107 ( .A(B[3]), .B(A[3]), .Z(n154) );
  IV U108 ( .A(n34), .Z(n140) );
  IVAP U109 ( .A(n140), .Z(n141) );
  IVDAP U110 ( .A(n6), .Y(n142), .Z(n143) );
  AN2P U111 ( .A(B[5]), .B(A[5]), .Z(n144) );
  MUX21HP U112 ( .A(n58), .B(n57), .S(n86), .Z(SUM[6]) );
  AN2P U113 ( .A(n149), .B(n150), .Z(n146) );
  EOP U114 ( .A(n165), .B(n164), .Z(n147) );
  IV U115 ( .A(n31), .Z(n27) );
  NR2P U116 ( .A(B[2]), .B(A[2]), .Z(n90) );
  AN2 U117 ( .A(A[8]), .B(B[8]), .Z(n148) );
  AN2 U118 ( .A(A[8]), .B(B[8]), .Z(n157) );
  IVP U119 ( .A(B[8]), .Z(n152) );
  ENP U120 ( .A(B[2]), .B(A[2]), .Z(SUM[2]) );
  IVDA U121 ( .A(A[4]), .Y(n149) );
  IV U122 ( .A(B[4]), .Z(n150) );
  AN2P U123 ( .A(A[7]), .B(B[7]), .Z(n50) );
  EOP U124 ( .A(n164), .B(n50), .Z(n159) );
  IV U125 ( .A(A[8]), .Z(n151) );
  ND2P U126 ( .A(n151), .B(n152), .Z(n156) );
  NR2P U127 ( .A(n8), .B(A[10]), .Z(n25) );
  ENP U128 ( .A(A[8]), .B(B[8]), .Z(n164) );
  ND2 U129 ( .A(n8), .B(A[10]), .Z(n26) );
  EOP U130 ( .A(A[7]), .B(B[7]), .Z(n51) );
  EOP U131 ( .A(B[5]), .B(A[5]), .Z(n162) );
  EOP U132 ( .A(B[9]), .B(A[9]), .Z(n33) );
  NR2P U133 ( .A(A[11]), .B(n143), .Z(n20) );
  EOP U134 ( .A(n19), .B(n26), .Z(n16) );
  EOP U135 ( .A(B[6]), .B(A[6]), .Z(n160) );
  EOP U136 ( .A(A[12]), .B(n143), .Z(n155) );
  EOP U137 ( .A(n8), .B(A[10]), .Z(n24) );
  EOP U138 ( .A(n25), .B(n19), .Z(n15) );
  MUX21L U139 ( .A(n148), .B(n156), .S(n165), .Z(n40) );
  IV U140 ( .A(n32), .Z(n28) );
  MUX21LP U141 ( .A(n60), .B(n59), .S(n86), .Z(n56) );
  MUX21LP U142 ( .A(n161), .B(n158), .S(n163), .Z(n63) );
  MUX21LP U143 ( .A(n161), .B(n158), .S(n144), .Z(n64) );
  IV U144 ( .A(n83), .Z(n80) );
  MUX21LP U145 ( .A(n71), .B(n72), .S(n84), .Z(SUM[5]) );
  ENP U146 ( .A(n79), .B(n162), .Z(n71) );
  MUX21LP U147 ( .A(n141), .B(n35), .S(n40), .Z(n31) );
  OR2P U148 ( .A(B[5]), .B(A[5]), .Z(n163) );
  OR2P U149 ( .A(B[6]), .B(A[6]), .Z(n158) );
  OR2P U150 ( .A(A[7]), .B(B[7]), .Z(n165) );
  IVP U151 ( .A(n56), .Z(n54) );
  MUX21L U152 ( .A(n63), .B(n64), .S(n83), .Z(n60) );
  MUX21L U153 ( .A(n63), .B(n64), .S(n146), .Z(n59) );
  MUX21L U154 ( .A(n18), .B(n17), .S(n31), .Z(n13) );
  MUX21L U155 ( .A(n18), .B(n17), .S(n32), .Z(n14) );
  EN U156 ( .A(n160), .B(n144), .Z(n62) );
  EN U157 ( .A(n163), .B(n160), .Z(n61) );
  MUX21L U158 ( .A(n11), .B(n12), .S(n56), .Z(SUM[11]) );
  MUX21L U159 ( .A(n16), .B(n15), .S(n31), .Z(n11) );
  MUX21L U160 ( .A(n16), .B(n15), .S(n32), .Z(n12) );
  MUX21L U161 ( .A(n61), .B(n62), .S(n83), .Z(n58) );
  MUX21L U162 ( .A(n61), .B(n62), .S(n146), .Z(n57) );
  IV U163 ( .A(n146), .Z(n79) );
  EO U164 ( .A(n90), .B(n154), .Z(SUM[3]) );
  MUX21L U165 ( .A(n23), .B(n22), .S(n54), .Z(SUM[10]) );
  EO U166 ( .A(n27), .B(n24), .Z(n22) );
  EO U167 ( .A(n28), .B(n24), .Z(n23) );
  EN U168 ( .A(A[4]), .B(B[4]), .Z(n81) );
  EO U169 ( .A(n40), .B(n33), .Z(n29) );
  EO U170 ( .A(n33), .B(n41), .Z(n30) );
  ND2 U171 ( .A(A[11]), .B(n143), .Z(n21) );
  EN U172 ( .A(A[11]), .B(n143), .Z(n19) );
  AN2P U173 ( .A(B[6]), .B(A[6]), .Z(n161) );
  OR2 U174 ( .A(A[12]), .B(A[13]), .Z(n166) );
  EOP U175 ( .A(n54), .B(n51), .Z(SUM[7]) );
  ND2 U176 ( .A(B[9]), .B(A[9]), .Z(n35) );
  ND2 U177 ( .A(B[3]), .B(A[3]), .Z(n89) );
  ND2 U178 ( .A(A[4]), .B(B[4]), .Z(n83) );
  IVAP U179 ( .A(n86), .Z(n84) );
endmodule


module prime_DW01_add_231 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n19, n20, n22, n24, n25, n26, n28, n30, n31, n32, n81, n82, n83, n84;

  ND2P U4 ( .A(B[12]), .B(B[13]), .Z(n7) );
  NR2 U7 ( .A(n12), .B(n11), .Z(n10) );
  EOP U10 ( .A(n20), .B(n1), .Z(SUM[5]) );
  ENP U20 ( .A(n2), .B(n25), .Z(SUM[4]) );
  MUX21LP U30 ( .A(n28), .B(n84), .S(n31), .Z(n26) );
  FA1A U37 ( .A(n32), .B(A[2]), .CI(B[2]), .CO(n31), .S(SUM[2]) );
  FA1A U38 ( .A(B[1]), .B(A[1]), .CI(n83), .CO(n32), .S(SUM[1]) );
  ND2 U46 ( .A(n10), .B(n13), .Z(n9) );
  NR2 U47 ( .A(n5), .B(n9), .Z(CO) );
  OR2P U48 ( .A(A[5]), .B(B[5]), .Z(n81) );
  IVA U49 ( .A(n24), .Z(n22) );
  OR2P U50 ( .A(A[4]), .B(B[4]), .Z(n82) );
  IV U51 ( .A(n30), .Z(n28) );
  OR2P U52 ( .A(B[0]), .B(A[0]), .Z(n83) );
  ND2 U53 ( .A(n81), .B(n19), .Z(n1) );
  ND2 U54 ( .A(B[11]), .B(B[10]), .Z(n8) );
  MUX21L U55 ( .A(n14), .B(n15), .S(n26), .Z(n13) );
  MUX21L U56 ( .A(n17), .B(n81), .S(n22), .Z(n15) );
  MUX21L U57 ( .A(n17), .B(n81), .S(n82), .Z(n14) );
  IVP U58 ( .A(n19), .Z(n17) );
  IV U59 ( .A(n26), .Z(n25) );
  ND2 U60 ( .A(n82), .B(n24), .Z(n2) );
  ND2 U61 ( .A(B[8]), .B(B[9]), .Z(n11) );
  MUX21L U62 ( .A(n22), .B(n82), .S(n25), .Z(n20) );
  ND2 U63 ( .A(B[7]), .B(B[6]), .Z(n12) );
  EN U64 ( .A(n3), .B(n31), .Z(SUM[3]) );
  ND2 U65 ( .A(n84), .B(n30), .Z(n3) );
  EN U66 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  OR2 U67 ( .A(A[3]), .B(B[3]), .Z(n84) );
  ND2 U68 ( .A(A[3]), .B(B[3]), .Z(n30) );
  ND2 U69 ( .A(n6), .B(B[14]), .Z(n5) );
  NR2P U70 ( .A(n8), .B(n7), .Z(n6) );
  ND2 U71 ( .A(A[5]), .B(B[5]), .Z(n19) );
  ND2 U72 ( .A(A[4]), .B(B[4]), .Z(n24) );
endmodule


module prime_DW01_add_224 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n14, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n36, n37, n38, n39,
         n40, n41, n45, n46, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n67, n68, n69, n70, n71, n72, n73,
         \A[0] , n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  AO6P U2 ( .A(n23), .B(n120), .C(n119), .Z(n9) );
  NR2 U10 ( .A(n21), .B(n19), .Z(n17) );
  NR2 U12 ( .A(A[11]), .B(B[11]), .Z(n19) );
  NR2 U14 ( .A(A[10]), .B(B[10]), .Z(n21) );
  AO7P U17 ( .A(n52), .B(n24), .C(n25), .Z(n23) );
  AO6P U19 ( .A(n39), .B(n26), .C(n27), .Z(n25) );
  NR2 U28 ( .A(n40), .B(n128), .Z(n31) );
  NR2 U54 ( .A(A[6]), .B(B[6]), .Z(n49) );
  AO6P U58 ( .A(n53), .B(n61), .C(n54), .Z(n52) );
  NR2 U59 ( .A(n58), .B(n55), .Z(n53) );
  NR2 U69 ( .A(A[4]), .B(B[4]), .Z(n58) );
  FA1A U79 ( .A(n130), .B(A[2]), .CI(B[2]), .CO(n64), .S(SUM[2]) );
  B5I U87 ( .A(n9), .Z(CO) );
  AN2 U88 ( .A(n18), .B(n14), .Z(n119) );
  AN2 U89 ( .A(n17), .B(n14), .Z(n120) );
  IVDA U90 ( .A(n50), .Y(n121), .Z(n122) );
  NR2P U91 ( .A(A[3]), .B(B[3]), .Z(n62) );
  AO7P U92 ( .A(n28), .B(n36), .C(n29), .Z(n27) );
  ND2P U93 ( .A(A[8]), .B(B[8]), .Z(n36) );
  ND2P U94 ( .A(n123), .B(n124), .Z(n125) );
  IVA U95 ( .A(A[8]), .Z(n123) );
  IVDA U96 ( .A(B[8]), .Y(n124) );
  IVAP U97 ( .A(n125), .Z(n128) );
  IV U98 ( .A(n72), .Z(n126) );
  NR2P U99 ( .A(n128), .B(n28), .Z(n26) );
  NR2 U100 ( .A(A[7]), .B(B[7]), .Z(n129) );
  NR2 U101 ( .A(A[7]), .B(B[7]), .Z(n127) );
  NR2P U102 ( .A(A[9]), .B(B[9]), .Z(n28) );
  AO7P U103 ( .A(n62), .B(n1), .C(n63), .Z(n61) );
  NR2P U104 ( .A(A[5]), .B(B[5]), .Z(n55) );
  IV U105 ( .A(n39), .Z(n41) );
  AO7P U106 ( .A(n129), .B(n50), .C(n45), .Z(n39) );
  AO7 U107 ( .A(n55), .B(n59), .C(n56), .Z(n54) );
  AO6P U108 ( .A(n51), .B(n31), .C(n32), .Z(n30) );
  EOP U109 ( .A(n30), .B(n2), .Z(SUM[9]) );
  IV U110 ( .A(n38), .Z(n40) );
  IV U111 ( .A(n61), .Z(n60) );
  ND2 U112 ( .A(n67), .B(n29), .Z(n2) );
  IV U113 ( .A(n52), .Z(n51) );
  EO U114 ( .A(n46), .B(n4), .Z(SUM[7]) );
  ND2 U115 ( .A(n69), .B(n45), .Z(n4) );
  EO U116 ( .A(n37), .B(n3), .Z(SUM[8]) );
  ND2 U117 ( .A(n68), .B(n36), .Z(n3) );
  AO6 U118 ( .A(n51), .B(n38), .C(n39), .Z(n37) );
  EN U119 ( .A(n57), .B(n6), .Z(SUM[5]) );
  IV U120 ( .A(n128), .Z(n68) );
  ND2 U121 ( .A(n71), .B(n56), .Z(n6) );
  IV U122 ( .A(n55), .Z(n71) );
  AN2P U123 ( .A(B[13]), .B(B[12]), .Z(n14) );
  NR2 U124 ( .A(n127), .B(n49), .Z(n38) );
  AO7 U125 ( .A(n19), .B(n22), .C(n20), .Z(n18) );
  ND2 U126 ( .A(A[11]), .B(B[11]), .Z(n20) );
  AO6 U127 ( .A(n51), .B(n70), .C(n121), .Z(n46) );
  EN U128 ( .A(n51), .B(n5), .Z(SUM[6]) );
  IV U129 ( .A(n49), .Z(n70) );
  ND2 U130 ( .A(n73), .B(n63), .Z(n8) );
  EO U131 ( .A(n7), .B(n60), .Z(SUM[4]) );
  ND2 U132 ( .A(n72), .B(n59), .Z(n7) );
  IVP U133 ( .A(n64), .Z(n1) );
  EN U134 ( .A(n8), .B(n64), .Z(SUM[3]) );
  OR2 U135 ( .A(B[1]), .B(A[1]), .Z(n130) );
  ND2 U136 ( .A(n70), .B(n122), .Z(n5) );
  IV U137 ( .A(n62), .Z(n73) );
  AO7 U138 ( .A(n60), .B(n126), .C(n59), .Z(n57) );
  IV U139 ( .A(n58), .Z(n72) );
  IV U140 ( .A(n28), .Z(n67) );
  IV U141 ( .A(n127), .Z(n69) );
  ND2 U142 ( .A(A[6]), .B(B[6]), .Z(n50) );
  ND2 U143 ( .A(A[3]), .B(B[3]), .Z(n63) );
  ND2 U144 ( .A(A[7]), .B(B[7]), .Z(n45) );
  ND2 U145 ( .A(A[10]), .B(B[10]), .Z(n22) );
  AO7 U146 ( .A(n41), .B(n128), .C(n36), .Z(n32) );
  ND2 U147 ( .A(n38), .B(n26), .Z(n24) );
  ND2 U148 ( .A(A[9]), .B(B[9]), .Z(n29) );
  ND2 U149 ( .A(A[5]), .B(B[5]), .Z(n56) );
  ND2 U150 ( .A(A[4]), .B(B[4]), .Z(n59) );
  EN U151 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
endmodule


module prime_DW01_add_223 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n9, n11, n15, n16, n17, n20, n21, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n41, n42,
         n45, n46, n47, n48, n49, \A[0] , \A[1] , n97, n98, n99, n100, n101,
         n102, n103, n104;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];

  MUX21LP U1 ( .A(n1), .B(n2), .S(n32), .Z(CO) );
  NR2 U10 ( .A(n104), .B(n11), .Z(n9) );
  NR2 U17 ( .A(A[8]), .B(B[8]), .Z(n15) );
  MUX21LP U37 ( .A(n36), .B(n35), .S(n45), .Z(n32) );
  MUX21LP U52 ( .A(n47), .B(n48), .S(n49), .Z(n45) );
  NR2 U57 ( .A(B[2]), .B(A[2]), .Z(n49) );
  EOP U62 ( .A(A[3]), .B(B[3]), .Z(n46) );
  EOP U63 ( .A(n17), .B(n98), .Z(SUM[8]) );
  ENP U64 ( .A(n46), .B(n49), .Z(SUM[3]) );
  EOP U65 ( .A(A[4]), .B(B[4]), .Z(n101) );
  NR2 U66 ( .A(A[6]), .B(B[6]), .Z(n97) );
  ND2P U67 ( .A(A[4]), .B(B[4]), .Z(n42) );
  EOP U68 ( .A(n37), .B(n42), .Z(n34) );
  EOP U69 ( .A(n45), .B(n101), .Z(SUM[4]) );
  MUX21LP U70 ( .A(n27), .B(n28), .S(n31), .Z(n25) );
  ND2P U71 ( .A(A[6]), .B(B[6]), .Z(n31) );
  MUX21L U72 ( .A(n27), .B(n28), .S(n30), .Z(n24) );
  NR2P U73 ( .A(A[7]), .B(B[7]), .Z(n27) );
  NR2P U74 ( .A(A[4]), .B(B[4]), .Z(n41) );
  NR2P U75 ( .A(A[6]), .B(B[6]), .Z(n30) );
  ENP U76 ( .A(n97), .B(n26), .Z(n100) );
  NR2P U77 ( .A(A[5]), .B(B[5]), .Z(n38) );
  IV U78 ( .A(n25), .Z(n21) );
  IV U79 ( .A(n24), .Z(n20) );
  MUX21L U80 ( .A(n4), .B(n3), .S(n25), .Z(n2) );
  EO U81 ( .A(A[8]), .B(B[8]), .Z(n98) );
  MUX21L U82 ( .A(n4), .B(n3), .S(n24), .Z(n1) );
  MUX21L U83 ( .A(n100), .B(n99), .S(n32), .Z(SUM[7]) );
  MUX21L U84 ( .A(n20), .B(n21), .S(n32), .Z(n17) );
  EN U85 ( .A(n26), .B(n31), .Z(n99) );
  ND2 U86 ( .A(A[7]), .B(B[7]), .Z(n28) );
  MUX21L U87 ( .A(n38), .B(n39), .S(n42), .Z(n36) );
  MUX21L U88 ( .A(n38), .B(n39), .S(n41), .Z(n35) );
  EO U89 ( .A(n32), .B(n29), .Z(SUM[6]) );
  EN U90 ( .A(A[6]), .B(B[6]), .Z(n29) );
  MUX21L U91 ( .A(n34), .B(n33), .S(n45), .Z(SUM[5]) );
  EO U92 ( .A(n41), .B(n37), .Z(n33) );
  EO U93 ( .A(A[5]), .B(B[5]), .Z(n37) );
  EN U94 ( .A(A[7]), .B(B[7]), .Z(n26) );
  ND2 U95 ( .A(B[9]), .B(B[10]), .Z(n11) );
  ND2 U96 ( .A(A[3]), .B(B[3]), .Z(n48) );
  ND2 U97 ( .A(n103), .B(B[13]), .Z(n102) );
  AN2P U98 ( .A(n9), .B(B[12]), .Z(n103) );
  EN U99 ( .A(B[2]), .B(A[2]), .Z(SUM[2]) );
  NR2P U100 ( .A(A[3]), .B(B[3]), .Z(n47) );
  NR2P U101 ( .A(n16), .B(n102), .Z(n4) );
  ND2 U102 ( .A(A[8]), .B(B[8]), .Z(n16) );
  ND2 U103 ( .A(A[5]), .B(B[5]), .Z(n39) );
  NR2P U104 ( .A(n15), .B(n102), .Z(n3) );
  IV U105 ( .A(B[11]), .Z(n104) );
endmodule


module prime_DW01_add_229 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n30, n31, n32,
         n34, n37, n38, n39, n40, n41, n42, n49, n50, n57, n58, n59, n60, n61,
         n62, n71, n74, n76, n78, n79, n80, n84, \B[1] , n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n150, n151,
         n152, n153, n154, n155, n156, n157, n159, n160;
  assign SUM[1] = \B[1] ;
  assign \B[1]  = B[1];

  ENP U2 ( .A(n2), .B(A[13]), .Z(SUM[13]) );
  MUX21LP U11 ( .A(n12), .B(n13), .S(n17), .Z(n9) );
  MUX21LP U12 ( .A(n160), .B(n13), .S(n18), .Z(n10) );
  EOP U17 ( .A(n19), .B(n16), .Z(n14) );
  EOP U18 ( .A(n20), .B(n16), .Z(n15) );
  MUX21LP U27 ( .A(n26), .B(n27), .S(n30), .Z(n23) );
  MUX21LP U28 ( .A(n26), .B(n27), .S(n31), .Z(n24) );
  MUX21LP U40 ( .A(n38), .B(n37), .S(n76), .Z(n34) );
  MUX21LP U55 ( .A(n49), .B(n50), .S(n74), .Z(SUM[7]) );
  ENP U56 ( .A(n57), .B(n139), .Z(n49) );
  ENP U57 ( .A(n58), .B(n139), .Z(n50) );
  MUX21LP U69 ( .A(n153), .B(n152), .S(n142), .Z(n61) );
  EOP U77 ( .A(n74), .B(n71), .Z(SUM[5]) );
  MUX21LP U86 ( .A(n78), .B(n79), .S(n80), .Z(n76) );
  NR2 U88 ( .A(A[4]), .B(B[4]), .Z(n78) );
  MUX21LP U91 ( .A(n141), .B(n137), .S(n138), .Z(n80) );
  ENP U104 ( .A(A[2]), .B(B[2]), .Z(SUM[2]) );
  OR2 U105 ( .A(B[3]), .B(A[3]), .Z(n137) );
  OR2P U106 ( .A(A[2]), .B(B[2]), .Z(n138) );
  EOP U107 ( .A(A[7]), .B(B[7]), .Z(n139) );
  EOP U108 ( .A(B[6]), .B(A[6]), .Z(n140) );
  AN2 U109 ( .A(B[3]), .B(A[3]), .Z(n141) );
  MUX21L U110 ( .A(n41), .B(n42), .S(n62), .Z(n38) );
  IV U111 ( .A(n62), .Z(n58) );
  MUX21LP U112 ( .A(n41), .B(n42), .S(n61), .Z(n37) );
  MUX21LP U113 ( .A(n59), .B(n60), .S(n74), .Z(SUM[6]) );
  ND2 U114 ( .A(B[10]), .B(A[10]), .Z(n27) );
  MUX21LP U115 ( .A(n3), .B(n4), .S(n148), .Z(SUM[12]) );
  ENP U116 ( .A(A[4]), .B(B[4]), .Z(n159) );
  EOP U117 ( .A(B[10]), .B(A[10]), .Z(n25) );
  EOP U118 ( .A(B[3]), .B(A[3]), .Z(n84) );
  OR2P U119 ( .A(n2), .B(A[13]), .Z(SUM[14]) );
  ENP U120 ( .A(A[9]), .B(B[9]), .Z(n147) );
  MUX21LP U121 ( .A(n39), .B(n40), .S(n62), .Z(n145) );
  MUX21LP U122 ( .A(n39), .B(n40), .S(n61), .Z(n146) );
  ENP U123 ( .A(n157), .B(n151), .Z(n39) );
  OR2 U124 ( .A(B[5]), .B(A[5]), .Z(n142) );
  OR2 U125 ( .A(B[5]), .B(A[5]), .Z(n143) );
  ENP U126 ( .A(n151), .B(n155), .Z(n40) );
  ND2 U127 ( .A(A[9]), .B(B[9]), .Z(n31) );
  IV U128 ( .A(n23), .Z(n19) );
  OR2 U129 ( .A(A[8]), .B(B[8]), .Z(n144) );
  OR2 U130 ( .A(A[8]), .B(B[8]), .Z(n150) );
  MUX21LP U131 ( .A(n156), .B(n144), .S(n157), .Z(n41) );
  MUX21LP U132 ( .A(n156), .B(n150), .S(n155), .Z(n42) );
  MUX21LP U133 ( .A(n14), .B(n15), .S(n148), .Z(SUM[11]) );
  EOP U134 ( .A(n25), .B(n30), .Z(n21) );
  EOP U135 ( .A(B[11]), .B(A[11]), .Z(n16) );
  NR2 U136 ( .A(A[11]), .B(B[11]), .Z(n17) );
  EOP U137 ( .A(B[8]), .B(A[8]), .Z(n151) );
  IVDAP U138 ( .A(n34), .Y(n32), .Z(n148) );
  EOP U139 ( .A(n17), .B(n11), .Z(n7) );
  NR2P U140 ( .A(A[12]), .B(B[12]), .Z(n160) );
  NR2P U141 ( .A(A[12]), .B(B[12]), .Z(n12) );
  ND2P U142 ( .A(A[12]), .B(B[12]), .Z(n13) );
  EOP U143 ( .A(n11), .B(n18), .Z(n8) );
  ENP U144 ( .A(A[12]), .B(B[12]), .Z(n11) );
  NR2P U145 ( .A(B[10]), .B(A[10]), .Z(n26) );
  EO U146 ( .A(n159), .B(n80), .Z(SUM[4]) );
  MUX21LP U147 ( .A(n153), .B(n152), .S(n154), .Z(n62) );
  MUX21H U148 ( .A(n145), .B(n146), .S(n76), .Z(SUM[8]) );
  EOP U149 ( .A(n34), .B(n147), .Z(SUM[9]) );
  MUX21LP U150 ( .A(n22), .B(n21), .S(n32), .Z(SUM[10]) );
  OR2P U151 ( .A(B[6]), .B(A[6]), .Z(n152) );
  OR2P U152 ( .A(A[7]), .B(B[7]), .Z(n157) );
  IV U153 ( .A(n61), .Z(n57) );
  EN U154 ( .A(n140), .B(n143), .Z(n59) );
  EN U155 ( .A(n140), .B(n154), .Z(n60) );
  EN U156 ( .A(A[6]), .B(A[5]), .Z(n71) );
  ND2 U157 ( .A(A[4]), .B(B[4]), .Z(n79) );
  MUX21L U158 ( .A(n8), .B(n7), .S(n23), .Z(n3) );
  MUX21L U159 ( .A(n8), .B(n7), .S(n24), .Z(n4) );
  AN2P U160 ( .A(B[6]), .B(A[6]), .Z(n153) );
  AN2P U161 ( .A(B[5]), .B(A[5]), .Z(n154) );
  AN2P U162 ( .A(A[7]), .B(B[7]), .Z(n155) );
  AN2P U163 ( .A(A[8]), .B(B[8]), .Z(n156) );
  EO U164 ( .A(n84), .B(n138), .Z(SUM[3]) );
  EO U165 ( .A(n25), .B(n31), .Z(n22) );
  IVA U166 ( .A(n24), .Z(n20) );
  MUX21L U167 ( .A(n10), .B(n9), .S(n24), .Z(n6) );
  MUX21L U168 ( .A(n10), .B(n9), .S(n23), .Z(n5) );
  NR2P U169 ( .A(A[9]), .B(B[9]), .Z(n30) );
  ND2 U170 ( .A(A[11]), .B(B[11]), .Z(n18) );
  MUX21L U171 ( .A(n5), .B(n6), .S(n34), .Z(n2) );
  IVAP U172 ( .A(n76), .Z(n74) );
endmodule


module prime_DW01_add_219 ( A, B, CI, SUM, CO );
  input [14:0] A;
  input [14:0] B;
  output [14:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n39, n40, n41, n46, n47, n48, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n60, n61, n62, n63, n64, n65, n66, n69, n71, n73, n75,
         \A[0] , n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n134;
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  NR2 U7 ( .A(n16), .B(n15), .Z(n14) );
  NR2 U12 ( .A(A[11]), .B(B[11]), .Z(n19) );
  NR2 U14 ( .A(A[10]), .B(B[10]), .Z(n21) );
  FA1A U81 ( .A(n134), .B(A[2]), .CI(B[2]), .CO(n66), .S(SUM[2]) );
  IVDA U89 ( .A(n60), .Y(n123), .Z(n124) );
  MUX21L U90 ( .A(n13), .B(n12), .S(n23), .Z(CO) );
  OR2 U91 ( .A(A[6]), .B(B[6]), .Z(n125) );
  ND2 U92 ( .A(A[8]), .B(B[8]), .Z(n127) );
  IVAP U93 ( .A(n130), .Z(n126) );
  MUX21LP U94 ( .A(n56), .B(n55), .S(n63), .Z(n130) );
  IV U95 ( .A(n63), .Z(n62) );
  ENP U96 ( .A(n8), .B(n66), .Z(SUM[3]) );
  ND2 U97 ( .A(A[3]), .B(B[3]), .Z(n65) );
  ND2 U98 ( .A(A[8]), .B(B[8]), .Z(n34) );
  MUX21L U99 ( .A(n28), .B(n29), .S(n33), .Z(n26) );
  IVDA U100 ( .A(n33), .Y(n129), .Z(n132) );
  IVDA U101 ( .A(n61), .Z(n128) );
  NR2P U102 ( .A(A[3]), .B(B[3]), .Z(n64) );
  NR2P U103 ( .A(A[9]), .B(B[9]), .Z(n28) );
  MUX21LP U104 ( .A(n46), .B(n47), .S(n51), .Z(n40) );
  MUX21LP U105 ( .A(n28), .B(n29), .S(n34), .Z(n27) );
  IVAP U106 ( .A(n54), .Z(n53) );
  MUX21LP U107 ( .A(n57), .B(n58), .S(n61), .Z(n56) );
  ND2P U108 ( .A(A[6]), .B(B[6]), .Z(n52) );
  MUX21LP U109 ( .A(n57), .B(n58), .S(n60), .Z(n55) );
  EOP U110 ( .A(n30), .B(n2), .Z(SUM[9]) );
  MUX21LP U111 ( .A(n56), .B(n55), .S(n63), .Z(n54) );
  NR2P U112 ( .A(A[7]), .B(B[7]), .Z(n46) );
  IV U113 ( .A(n52), .Z(n50) );
  EOP U114 ( .A(n131), .B(n6), .Z(SUM[5]) );
  MUX21H U115 ( .A(n124), .B(n128), .S(n62), .Z(n131) );
  MUX21LP U116 ( .A(n65), .B(n64), .S(n66), .Z(n63) );
  NR2P U117 ( .A(A[8]), .B(B[8]), .Z(n33) );
  MUX21L U118 ( .A(n127), .B(n132), .S(n40), .Z(n31) );
  MUX21L U119 ( .A(n127), .B(n132), .S(n41), .Z(n32) );
  IVP U120 ( .A(n46), .Z(n71) );
  EO U121 ( .A(n39), .B(n3), .Z(SUM[8]) );
  ND2 U122 ( .A(n129), .B(n127), .Z(n3) );
  MUX21L U123 ( .A(n41), .B(n40), .S(n53), .Z(n39) );
  MUX21L U124 ( .A(n46), .B(n47), .S(n52), .Z(n41) );
  ND2 U125 ( .A(n69), .B(n29), .Z(n2) );
  MUX21L U126 ( .A(n32), .B(n31), .S(n126), .Z(n30) );
  IV U127 ( .A(n28), .Z(n69) );
  ND2 U128 ( .A(A[7]), .B(B[7]), .Z(n47) );
  EN U129 ( .A(n53), .B(n5), .Z(SUM[6]) );
  ND2 U130 ( .A(n125), .B(n52), .Z(n5) );
  MUX21L U131 ( .A(n24), .B(n25), .S(n130), .Z(n23) );
  MUX21L U132 ( .A(n27), .B(n26), .S(n40), .Z(n24) );
  MUX21L U133 ( .A(n27), .B(n26), .S(n41), .Z(n25) );
  ND2 U134 ( .A(A[9]), .B(B[9]), .Z(n29) );
  ND2 U135 ( .A(n17), .B(n14), .Z(n12) );
  MUX21L U136 ( .A(n19), .B(n20), .S(n21), .Z(n17) );
  ND2 U137 ( .A(n18), .B(n14), .Z(n13) );
  MUX21L U138 ( .A(n19), .B(n20), .S(n22), .Z(n18) );
  ND2 U139 ( .A(A[10]), .B(B[10]), .Z(n22) );
  ND2 U140 ( .A(n73), .B(n58), .Z(n6) );
  IV U141 ( .A(n57), .Z(n73) );
  ND2 U142 ( .A(A[11]), .B(B[11]), .Z(n20) );
  ND2 U143 ( .A(n123), .B(n128), .Z(n7) );
  IVDA U144 ( .A(B[14]), .Y(n15) );
  EO U145 ( .A(n7), .B(n62), .Z(SUM[4]) );
  EO U146 ( .A(n48), .B(n4), .Z(SUM[7]) );
  ND2 U147 ( .A(n71), .B(n47), .Z(n4) );
  MUX21L U148 ( .A(n50), .B(n125), .S(n53), .Z(n48) );
  OR2 U149 ( .A(B[1]), .B(A[1]), .Z(n134) );
  EN U150 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  ND2 U151 ( .A(n75), .B(n65), .Z(n8) );
  IV U152 ( .A(n64), .Z(n75) );
  NR2P U153 ( .A(A[5]), .B(B[5]), .Z(n57) );
  ND2 U154 ( .A(A[5]), .B(B[5]), .Z(n58) );
  NR2P U155 ( .A(A[6]), .B(B[6]), .Z(n51) );
  ND2 U156 ( .A(B[13]), .B(B[12]), .Z(n16) );
  ND2 U157 ( .A(A[4]), .B(B[4]), .Z(n61) );
  NR2P U158 ( .A(A[4]), .B(B[4]), .Z(n60) );
endmodule


module prime_DW01_sub_8 ( A, B, CI, DIFF, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] DIFF;
  input CI;
  output CO;
  wire   n2, n6, n7, n12, n13, n14, n16, n17, n18, n19, n20, n26, n27, n37,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n67, n68, n69,
         n70, n72, n75, n76, n77, n78, n79, n81, n82, n85, n87, n88, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n162, n163, n164, n165, n167, n168, n169, n170, n171, n172, n173,
         n174, n176;
  assign n14 = B[9];
  assign n20 = B[8];
  assign n87 = B[2];

  EOP U4 ( .A(n12), .B(A[13]), .Z(n6) );
  MUX21LP U16 ( .A(n17), .B(n16), .S(n2), .Z(DIFF[11]) );
  MUX21LP U45 ( .A(n43), .B(n44), .S(n72), .Z(n2) );
  NR2 U55 ( .A(n169), .B(A[8]), .Z(n50) );
  MUX21LP U57 ( .A(n53), .B(n52), .S(n70), .Z(DIFF[7]) );
  EOP U58 ( .A(n57), .B(n54), .Z(n52) );
  EOP U59 ( .A(n58), .B(n54), .Z(n53) );
  MUX21LP U63 ( .A(n60), .B(n59), .S(n70), .Z(DIFF[6]) );
  MUX21LP U68 ( .A(n64), .B(n65), .S(n68), .Z(n61) );
  MUX21LP U69 ( .A(n64), .B(n65), .S(n69), .Z(n62) );
  ND2P U77 ( .A(n172), .B(A[5]), .Z(n69) );
  MUX21LP U81 ( .A(n76), .B(n75), .S(n85), .Z(n72) );
  NR2 U100 ( .A(n176), .B(n149), .Z(n88) );
  MUX21L U118 ( .A(n78), .B(n79), .S(n82), .Z(n76) );
  B3I U119 ( .A(B[0]), .Z1(n149), .Z2(n150) );
  EOP U120 ( .A(n18), .B(n168), .Z(n151) );
  EOP U121 ( .A(n165), .B(n159), .Z(n152) );
  NR2P U122 ( .A(n26), .B(n169), .Z(n18) );
  NR2P U123 ( .A(n27), .B(n169), .Z(n19) );
  MUX21LP U124 ( .A(n156), .B(n151), .S(n153), .Z(DIFF[12]) );
  NR2P U125 ( .A(n170), .B(A[7]), .Z(n55) );
  NR2P U126 ( .A(n171), .B(A[6]), .Z(n64) );
  ENP U127 ( .A(n176), .B(n149), .Z(DIFF[1]) );
  MUX21L U128 ( .A(n50), .B(n51), .S(n56), .Z(n48) );
  EOP U129 ( .A(n55), .B(n49), .Z(n45) );
  ENP U130 ( .A(n169), .B(A[8]), .Z(n49) );
  ND2P U131 ( .A(A[4]), .B(n173), .Z(n79) );
  ENP U132 ( .A(A[4]), .B(n173), .Z(n77) );
  EOP U133 ( .A(n170), .B(A[7]), .Z(n54) );
  AN2P U134 ( .A(B[3]), .B(n149), .Z(n81) );
  AN2P U135 ( .A(n176), .B(B[4]), .Z(n78) );
  MUX21LP U136 ( .A(n43), .B(n44), .S(n72), .Z(n153) );
  OR2P U137 ( .A(n154), .B(n149), .Z(n85) );
  ND2 U138 ( .A(B[1]), .B(n87), .Z(n154) );
  MUX21LP U139 ( .A(n48), .B(n47), .S(n61), .Z(n43) );
  EOP U140 ( .A(n13), .B(A[13]), .Z(n7) );
  IV U141 ( .A(B[10]), .Z(n167) );
  IVP U142 ( .A(B[3]), .Z(n174) );
  IV U143 ( .A(B[1]), .Z(n176) );
  B5I U144 ( .A(B[7]), .Z(n170) );
  ENP U145 ( .A(n88), .B(n87), .Z(DIFF[2]) );
  EN U146 ( .A(n77), .B(n81), .Z(n163) );
  MUX21LP U147 ( .A(n155), .B(n152), .S(n2), .Z(DIFF[10]) );
  MUX21L U148 ( .A(n7), .B(n6), .S(n153), .Z(DIFF[13]) );
  MUX21L U149 ( .A(n48), .B(n47), .S(n62), .Z(n44) );
  ND2P U150 ( .A(n174), .B(A[3]), .Z(n82) );
  NR2P U151 ( .A(n172), .B(A[5]), .Z(n68) );
  IVAP U152 ( .A(n72), .Z(n70) );
  EO U153 ( .A(n159), .B(n164), .Z(n155) );
  EO U154 ( .A(n19), .B(n168), .Z(n156) );
  OR2P U155 ( .A(n167), .B(A[10]), .Z(n157) );
  MUX21L U156 ( .A(n50), .B(n51), .S(n55), .Z(n47) );
  IV U157 ( .A(n62), .Z(n58) );
  MUX21L U158 ( .A(n158), .B(n157), .S(n164), .Z(n27) );
  MUX21L U159 ( .A(n158), .B(n157), .S(n165), .Z(n26) );
  ND2 U160 ( .A(n170), .B(A[7]), .Z(n56) );
  ND2 U161 ( .A(n169), .B(A[8]), .Z(n51) );
  EO U162 ( .A(n171), .B(A[6]), .Z(n63) );
  MUX21L U163 ( .A(n41), .B(n42), .S(n72), .Z(DIFF[8]) );
  MUX21L U164 ( .A(n46), .B(n45), .S(n61), .Z(n41) );
  MUX21L U165 ( .A(n46), .B(n45), .S(n62), .Z(n42) );
  EO U166 ( .A(n49), .B(n56), .Z(n46) );
  AN2P U167 ( .A(n167), .B(A[10]), .Z(n158) );
  EN U168 ( .A(n167), .B(A[10]), .Z(n159) );
  EO U169 ( .A(n85), .B(n160), .Z(DIFF[3]) );
  EO U170 ( .A(n174), .B(n150), .Z(n160) );
  EOP U171 ( .A(n70), .B(n67), .Z(DIFF[5]) );
  EO U172 ( .A(n172), .B(A[5]), .Z(n67) );
  EOP U173 ( .A(n2), .B(n37), .Z(DIFF[9]) );
  EO U174 ( .A(n168), .B(A[9]), .Z(n37) );
  MUX21L U175 ( .A(n162), .B(n163), .S(n85), .Z(DIFF[4]) );
  EN U176 ( .A(n77), .B(n82), .Z(n162) );
  EO U177 ( .A(n27), .B(n20), .Z(n17) );
  EO U178 ( .A(n26), .B(n20), .Z(n16) );
  MUX21L U179 ( .A(n78), .B(n79), .S(n81), .Z(n75) );
  AN2P U180 ( .A(n168), .B(A[9]), .Z(n164) );
  OR2 U181 ( .A(n168), .B(A[9]), .Z(n165) );
  IV U182 ( .A(B[5]), .Z(n172) );
  IV U183 ( .A(B[4]), .Z(n173) );
  EO U184 ( .A(n63), .B(n69), .Z(n60) );
  EO U185 ( .A(n68), .B(n63), .Z(n59) );
  IVP U186 ( .A(n61), .Z(n57) );
  ND2 U187 ( .A(n19), .B(n14), .Z(n13) );
  ND2 U188 ( .A(n18), .B(n14), .Z(n12) );
  ND2 U189 ( .A(n171), .B(A[6]), .Z(n65) );
  IVA U190 ( .A(n14), .Z(n168) );
  IVA U191 ( .A(n20), .Z(n169) );
  IVA U192 ( .A(B[6]), .Z(n171) );
  IV U193 ( .A(n149), .Z(DIFF[0]) );
endmodule


module prime_DW01_add_240 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n3, n4, n5, n6, n8, n11, n12, n13, n14, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n48, n49, n50, n51, n53,
         n56, n57, n58, n59, n60, n62, n63, n66, n68, n69, n70, \B[0] , \B[1] ,
         n117, n119, n120, n122, n123, n124, n125, n126, n127;
  assign n8 = B[10];
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];
  assign SUM[1] = \B[1] ;
  assign \B[1]  = B[1];

  NR2 U7 ( .A(n13), .B(n123), .Z(n5) );
  NR2 U8 ( .A(n14), .B(n123), .Z(n6) );
  NR2 U23 ( .A(A[10]), .B(n123), .Z(n19) );
  MUX21LP U26 ( .A(n24), .B(n25), .S(n53), .Z(n21) );
  EOP U32 ( .A(n30), .B(n37), .Z(n27) );
  MUX21LP U34 ( .A(n31), .B(n32), .S(n37), .Z(n29) );
  NR2 U36 ( .A(A[9]), .B(n125), .Z(n31) );
  MUX21LP U38 ( .A(n34), .B(n33), .S(n51), .Z(SUM[8]) );
  EOP U39 ( .A(n38), .B(n35), .Z(n33) );
  EOP U40 ( .A(n39), .B(n35), .Z(n34) );
  NR2 U42 ( .A(A[8]), .B(B[8]), .Z(n36) );
  MUX21LP U44 ( .A(n41), .B(n40), .S(n51), .Z(SUM[7]) );
  MUX21LP U49 ( .A(n45), .B(n46), .S(n49), .Z(n42) );
  MUX21LP U62 ( .A(n57), .B(n56), .S(n66), .Z(n53) );
  MUX21LP U77 ( .A(n68), .B(n69), .S(n70), .Z(n66) );
  NR2 U79 ( .A(A[3]), .B(B[3]), .Z(n68) );
  MUX21L U86 ( .A(n6), .B(n5), .S(n21), .Z(SUM[13]) );
  ND2P U87 ( .A(A[6]), .B(B[6]), .Z(n50) );
  NR2P U88 ( .A(A[4]), .B(B[4]), .Z(n62) );
  EOP U89 ( .A(A[7]), .B(B[7]), .Z(n44) );
  NR2P U90 ( .A(A[7]), .B(B[7]), .Z(n45) );
  NR2 U91 ( .A(A[5]), .B(B[5]), .Z(n59) );
  EOP U92 ( .A(A[6]), .B(B[6]), .Z(n48) );
  ENP U93 ( .A(A[5]), .B(B[5]), .Z(n58) );
  EOP U94 ( .A(A[4]), .B(B[4]), .Z(n117) );
  ENP U95 ( .A(n62), .B(n58), .Z(n120) );
  ENP U96 ( .A(n58), .B(n63), .Z(n119) );
  EOP U97 ( .A(n66), .B(n117), .Z(SUM[4]) );
  EOP U98 ( .A(n49), .B(n44), .Z(n40) );
  NR2P U99 ( .A(A[6]), .B(B[6]), .Z(n49) );
  ENP U100 ( .A(A[2]), .B(B[2]), .Z(SUM[2]) );
  ENP U101 ( .A(A[3]), .B(B[3]), .Z(n122) );
  IVA U102 ( .A(n53), .Z(n51) );
  NR2P U103 ( .A(A[2]), .B(B[2]), .Z(n70) );
  IV U104 ( .A(n42), .Z(n38) );
  EOP U105 ( .A(n36), .B(n30), .Z(n26) );
  MUX21LP U106 ( .A(n45), .B(n46), .S(n50), .Z(n43) );
  MUX21LP U107 ( .A(n31), .B(n32), .S(n36), .Z(n28) );
  IVAP U108 ( .A(n126), .Z(n125) );
  IVP U109 ( .A(n43), .Z(n39) );
  MUX21L U110 ( .A(n12), .B(n11), .S(n21), .Z(SUM[11]) );
  EO U111 ( .A(n20), .B(n127), .Z(n12) );
  EO U112 ( .A(n19), .B(n127), .Z(n11) );
  MUX21H U113 ( .A(n4), .B(n3), .S(n21), .Z(SUM[12]) );
  EN U114 ( .A(n14), .B(n123), .Z(n4) );
  EO U115 ( .A(n44), .B(n50), .Z(n41) );
  ND2 U116 ( .A(A[9]), .B(n125), .Z(n32) );
  EN U117 ( .A(n13), .B(n123), .Z(n3) );
  EN U118 ( .A(A[9]), .B(n125), .Z(n30) );
  ND2 U119 ( .A(n20), .B(n127), .Z(n14) );
  ND2 U120 ( .A(n19), .B(n127), .Z(n13) );
  EOP U121 ( .A(n21), .B(n18), .Z(SUM[10]) );
  EO U122 ( .A(A[10]), .B(n123), .Z(n18) );
  MUX21L U123 ( .A(n29), .B(n28), .S(n42), .Z(n24) );
  MUX21L U124 ( .A(n29), .B(n28), .S(n43), .Z(n25) );
  MUX21L U125 ( .A(n119), .B(n120), .S(n66), .Z(SUM[5]) );
  EOP U126 ( .A(n51), .B(n48), .Z(SUM[6]) );
  EO U127 ( .A(n122), .B(n70), .Z(SUM[3]) );
  ND2 U128 ( .A(A[4]), .B(B[4]), .Z(n63) );
  EO U129 ( .A(A[8]), .B(B[8]), .Z(n35) );
  ND2 U130 ( .A(A[8]), .B(B[8]), .Z(n37) );
  MUX21L U131 ( .A(n22), .B(n23), .S(n53), .Z(SUM[9]) );
  MUX21L U132 ( .A(n27), .B(n26), .S(n42), .Z(n22) );
  MUX21L U133 ( .A(n27), .B(n26), .S(n43), .Z(n23) );
  ND2 U134 ( .A(A[10]), .B(n123), .Z(n20) );
  ND2 U135 ( .A(A[7]), .B(B[7]), .Z(n46) );
  ND2 U136 ( .A(A[3]), .B(B[3]), .Z(n69) );
  MUX21L U137 ( .A(n59), .B(n60), .S(n63), .Z(n57) );
  MUX21L U138 ( .A(n59), .B(n60), .S(n62), .Z(n56) );
  ND2 U139 ( .A(A[5]), .B(B[5]), .Z(n60) );
  IVA U140 ( .A(n124), .Z(n123) );
  IV U141 ( .A(n8), .Z(n124) );
  IVA U142 ( .A(B[9]), .Z(n126) );
  IVA U143 ( .A(n125), .Z(n127) );
endmodule


module prime_DW01_add_215 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n8, n13, n14, n15, n16, n17, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n51, n52, n54, n57,
         n58, n59, n60, n61, n63, n64, n67, n69, n70, n71, \B[1] , n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n132, n133, n134, n136, n137, n138;
  assign n8 = B[11];
  assign SUM[1] = \B[1] ;
  assign \B[1]  = B[1];

  MUX21LP U1 ( .A(n6), .B(n5), .S(n127), .Z(SUM[13]) );
  MUX21LP U2 ( .A(n130), .B(n119), .S(n127), .Z(SUM[12]) );
  NR2 U7 ( .A(n13), .B(n137), .Z(n5) );
  NR2 U8 ( .A(n14), .B(n137), .Z(n6) );
  MUX21LP U16 ( .A(n16), .B(n17), .S(n20), .Z(n13) );
  MUX21LP U17 ( .A(n16), .B(n17), .S(n21), .Z(n14) );
  EOP U18 ( .A(n137), .B(A[11]), .Z(n15) );
  NR2 U24 ( .A(A[10]), .B(B[10]), .Z(n20) );
  MUX21LP U34 ( .A(n32), .B(n33), .S(n37), .Z(n29) );
  MUX21LP U35 ( .A(n32), .B(n33), .S(n38), .Z(n30) );
  MUX21LP U39 ( .A(n35), .B(n34), .S(n52), .Z(SUM[8]) );
  EOP U40 ( .A(n120), .B(n36), .Z(n34) );
  EOP U41 ( .A(n40), .B(n36), .Z(n35) );
  MUX21LP U50 ( .A(n46), .B(n47), .S(n50), .Z(n43) );
  MUX21LP U51 ( .A(n46), .B(n47), .S(n51), .Z(n44) );
  ND2P U59 ( .A(A[6]), .B(B[6]), .Z(n51) );
  MUX21LP U63 ( .A(n58), .B(n57), .S(n67), .Z(n54) );
  MUX21LP U78 ( .A(n69), .B(n70), .S(n71), .Z(n67) );
  NR2 U80 ( .A(A[3]), .B(B[3]), .Z(n69) );
  MUX21L U87 ( .A(n25), .B(n26), .S(n54), .Z(n22) );
  MUX21L U88 ( .A(n28), .B(n27), .S(n122), .Z(n23) );
  IVDA U89 ( .A(A[2]), .Z(n118) );
  EOP U90 ( .A(n13), .B(n137), .Z(n119) );
  EN U91 ( .A(B[3]), .B(A[3]), .Z(n136) );
  IVDA U92 ( .A(B[2]), .Z(n121) );
  IVDA U93 ( .A(n43), .Y(n120), .Z(n122) );
  EOP U94 ( .A(A[6]), .B(B[6]), .Z(n49) );
  NR2P U95 ( .A(A[9]), .B(B[9]), .Z(n32) );
  MUX21LP U96 ( .A(n60), .B(n61), .S(n63), .Z(n57) );
  NR2 U97 ( .A(B[5]), .B(A[5]), .Z(n60) );
  NR2 U98 ( .A(n121), .B(A[2]), .Z(n123) );
  MUX21LP U99 ( .A(n58), .B(n57), .S(n67), .Z(n124) );
  IVDA U100 ( .A(n67), .Z(n126) );
  EOP U101 ( .A(B[7]), .B(A[7]), .Z(n45) );
  MUX21L U102 ( .A(n30), .B(n29), .S(n43), .Z(n125) );
  MUX21L U103 ( .A(n30), .B(n29), .S(n43), .Z(n25) );
  EO U104 ( .A(n50), .B(n45), .Z(n41) );
  IVAP U105 ( .A(n124), .Z(n52) );
  EOP U106 ( .A(A[10]), .B(B[10]), .Z(n19) );
  NR2 U107 ( .A(n137), .B(A[11]), .Z(n16) );
  NR2 U108 ( .A(A[4]), .B(B[4]), .Z(n63) );
  NR2P U109 ( .A(B[7]), .B(A[7]), .Z(n46) );
  ENP U110 ( .A(n121), .B(n118), .Z(SUM[2]) );
  EOP U111 ( .A(n136), .B(n123), .Z(SUM[3]) );
  NR2P U112 ( .A(A[8]), .B(B[8]), .Z(n37) );
  EOP U113 ( .A(n37), .B(n31), .Z(n27) );
  EOP U114 ( .A(A[4]), .B(B[4]), .Z(n134) );
  IVAP U115 ( .A(n138), .Z(n137) );
  ENP U116 ( .A(B[5]), .B(A[5]), .Z(n59) );
  MUX21LP U117 ( .A(n23), .B(n24), .S(n124), .Z(SUM[9]) );
  EOP U118 ( .A(n67), .B(n134), .Z(SUM[4]) );
  MUX21LP U119 ( .A(n125), .B(n26), .S(n54), .Z(n127) );
  MUX21LP U120 ( .A(n30), .B(n29), .S(n44), .Z(n26) );
  MUX21LP U121 ( .A(n128), .B(n129), .S(n22), .Z(SUM[11]) );
  EOP U122 ( .A(n31), .B(n38), .Z(n28) );
  MUX21LP U123 ( .A(n132), .B(n133), .S(n126), .Z(SUM[5]) );
  ENP U124 ( .A(n63), .B(n59), .Z(n133) );
  MUX21LP U125 ( .A(n42), .B(n41), .S(n52), .Z(SUM[7]) );
  EO U126 ( .A(n15), .B(n21), .Z(n128) );
  EO U127 ( .A(n20), .B(n15), .Z(n129) );
  EO U128 ( .A(n14), .B(n137), .Z(n130) );
  MUX21L U129 ( .A(n28), .B(n27), .S(n44), .Z(n24) );
  IV U130 ( .A(n44), .Z(n40) );
  EOP U131 ( .A(n22), .B(n19), .Z(SUM[10]) );
  EN U132 ( .A(n59), .B(n64), .Z(n132) );
  MUX21L U133 ( .A(n60), .B(n61), .S(n64), .Z(n58) );
  ND2 U134 ( .A(B[5]), .B(A[5]), .Z(n61) );
  ND2 U135 ( .A(B[7]), .B(A[7]), .Z(n47) );
  ND2 U136 ( .A(A[8]), .B(B[8]), .Z(n38) );
  EO U137 ( .A(A[8]), .B(B[8]), .Z(n36) );
  EO U138 ( .A(n45), .B(n51), .Z(n42) );
  ND2 U139 ( .A(A[9]), .B(B[9]), .Z(n33) );
  EN U140 ( .A(A[9]), .B(B[9]), .Z(n31) );
  EOP U141 ( .A(n52), .B(n49), .Z(SUM[6]) );
  ND2 U142 ( .A(A[4]), .B(B[4]), .Z(n64) );
  ND2 U143 ( .A(n137), .B(A[11]), .Z(n17) );
  ND2 U144 ( .A(A[10]), .B(B[10]), .Z(n21) );
  ND2 U145 ( .A(A[3]), .B(B[3]), .Z(n70) );
  NR2P U146 ( .A(A[6]), .B(B[6]), .Z(n50) );
  NR2P U147 ( .A(B[2]), .B(A[2]), .Z(n71) );
  IV U148 ( .A(n8), .Z(n138) );
endmodule


module prime_DW01_add_217 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n5, n6, n8, n11, n12, n13, n14, n15, n16, n17, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n51,
         n52, n54, n57, n58, n59, n61, n63, n64, n67, n69, n70, n71, \B[0] ,
         n118, n119, n120, n121, n122, n123, n125, n126, n128, n129, n130,
         n131;
  assign n8 = B[10];
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  MUX21LP U2 ( .A(n123), .B(n118), .S(n22), .Z(SUM[11]) );
  NR2 U7 ( .A(n13), .B(n130), .Z(n5) );
  NR2 U8 ( .A(n14), .B(n130), .Z(n6) );
  NR2 U19 ( .A(n130), .B(A[10]), .Z(n16) );
  NR2 U24 ( .A(A[9]), .B(B[9]), .Z(n20) );
  MUX21LP U27 ( .A(n25), .B(n26), .S(n54), .Z(n22) );
  NR2 U37 ( .A(A[8]), .B(B[8]), .Z(n32) );
  EOP U40 ( .A(n39), .B(n36), .Z(n34) );
  EOP U41 ( .A(n40), .B(n36), .Z(n35) );
  NR2 U43 ( .A(A[7]), .B(B[7]), .Z(n37) );
  MUX21LP U51 ( .A(n46), .B(n47), .S(n51), .Z(n44) );
  MUX21LP U63 ( .A(n58), .B(n57), .S(n67), .Z(n54) );
  MUX21LP U78 ( .A(n69), .B(n70), .S(n71), .Z(n67) );
  EOP U87 ( .A(n13), .B(n130), .Z(n118) );
  NR2P U88 ( .A(B[4]), .B(A[4]), .Z(n119) );
  NR2 U89 ( .A(B[1]), .B(A[1]), .Z(n120) );
  ENP U90 ( .A(A[1]), .B(B[1]), .Z(SUM[1]) );
  EOP U91 ( .A(B[6]), .B(A[6]), .Z(n45) );
  EO U92 ( .A(A[5]), .B(B[5]), .Z(n49) );
  IVDA U93 ( .A(n51), .Z(n122) );
  MUX21LP U94 ( .A(n119), .B(n61), .S(n63), .Z(n57) );
  MUX21LP U95 ( .A(n119), .B(n61), .S(n64), .Z(n58) );
  ENP U96 ( .A(n121), .B(n49), .Z(SUM[5]) );
  EOP U97 ( .A(n130), .B(A[10]), .Z(n15) );
  MUX21LP U98 ( .A(n125), .B(n126), .S(n67), .Z(SUM[4]) );
  NR2 U99 ( .A(A[3]), .B(B[3]), .Z(n63) );
  NR2P U100 ( .A(B[6]), .B(A[6]), .Z(n46) );
  MUX21LP U101 ( .A(n58), .B(n57), .S(n67), .Z(n121) );
  IVAP U102 ( .A(n121), .Z(n52) );
  MUX21LP U103 ( .A(n35), .B(n34), .S(n52), .Z(SUM[7]) );
  NR2P U104 ( .A(A[2]), .B(B[2]), .Z(n69) );
  ENP U105 ( .A(B[4]), .B(A[4]), .Z(n59) );
  EOP U106 ( .A(A[3]), .B(B[3]), .Z(n129) );
  ENP U107 ( .A(A[2]), .B(B[2]), .Z(n128) );
  ENP U108 ( .A(n63), .B(n59), .Z(n126) );
  NR2P U109 ( .A(A[5]), .B(B[5]), .Z(n50) );
  NR2P U110 ( .A(B[1]), .B(A[1]), .Z(n71) );
  EOP U111 ( .A(n128), .B(n120), .Z(SUM[2]) );
  IV U112 ( .A(n44), .Z(n40) );
  MUX21LP U113 ( .A(n46), .B(n47), .S(n50), .Z(n43) );
  MUX21LP U114 ( .A(n16), .B(n17), .S(n20), .Z(n13) );
  IVP U115 ( .A(n43), .Z(n39) );
  MUX21L U116 ( .A(n6), .B(n5), .S(n22), .Z(SUM[12]) );
  EO U117 ( .A(n14), .B(n130), .Z(n123) );
  MUX21L U118 ( .A(n30), .B(n29), .S(n44), .Z(n26) );
  MUX21L U119 ( .A(n30), .B(n29), .S(n43), .Z(n25) );
  MUX21L U120 ( .A(n32), .B(n33), .S(n38), .Z(n30) );
  MUX21L U121 ( .A(n23), .B(n24), .S(n54), .Z(SUM[8]) );
  MUX21L U122 ( .A(n28), .B(n27), .S(n44), .Z(n24) );
  MUX21L U123 ( .A(n28), .B(n27), .S(n43), .Z(n23) );
  EO U124 ( .A(n31), .B(n38), .Z(n28) );
  ND2 U125 ( .A(A[5]), .B(B[5]), .Z(n51) );
  MUX21L U126 ( .A(n32), .B(n33), .S(n37), .Z(n29) );
  MUX21L U127 ( .A(n16), .B(n17), .S(n21), .Z(n14) );
  EO U128 ( .A(n37), .B(n31), .Z(n27) );
  EOP U129 ( .A(n22), .B(n19), .Z(SUM[9]) );
  EO U130 ( .A(A[9]), .B(B[9]), .Z(n19) );
  MUX21L U131 ( .A(n12), .B(n11), .S(n22), .Z(SUM[10]) );
  EO U132 ( .A(n15), .B(n21), .Z(n12) );
  EO U133 ( .A(n20), .B(n15), .Z(n11) );
  ND2 U134 ( .A(B[4]), .B(A[4]), .Z(n61) );
  EN U135 ( .A(n59), .B(n64), .Z(n125) );
  EO U136 ( .A(A[7]), .B(B[7]), .Z(n36) );
  MUX21L U137 ( .A(n42), .B(n41), .S(n52), .Z(SUM[6]) );
  EO U138 ( .A(n45), .B(n122), .Z(n42) );
  EO U139 ( .A(n50), .B(n45), .Z(n41) );
  ND2 U140 ( .A(B[6]), .B(A[6]), .Z(n47) );
  ND2 U141 ( .A(A[7]), .B(B[7]), .Z(n38) );
  ND2 U142 ( .A(A[8]), .B(B[8]), .Z(n33) );
  EN U143 ( .A(A[8]), .B(B[8]), .Z(n31) );
  EO U144 ( .A(n67), .B(n129), .Z(SUM[3]) );
  ND2 U145 ( .A(A[2]), .B(B[2]), .Z(n70) );
  ND2 U146 ( .A(n130), .B(A[10]), .Z(n17) );
  ND2 U147 ( .A(A[9]), .B(B[9]), .Z(n21) );
  ND2 U148 ( .A(A[3]), .B(B[3]), .Z(n64) );
  IVA U149 ( .A(n131), .Z(n130) );
  IV U150 ( .A(n8), .Z(n131) );
endmodule


module prime_add_0_root_add_212_I6_DP_OP_297_0_0 ( I1, I2, I3, I4, I5, I6, O2
 );
  input [1:0] I1;
  input [11:0] I2;
  input [9:0] I3;
  input [7:0] I4;
  input [5:0] I5;
  input [3:0] I6;
  output [13:0] O2;
  wire   n62, n67, n70, n71, n72, n73, n74, n76, n77, n80, n82, n83, n84, n98,
         n99, n113, n115, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n158, n194, n195, n196, n197, n198, n199, n200, n201, n206, n207,
         n209, n210, n211, n212, n213;
  assign O2[5] = n158;
  assign n194 = I2[2];
  assign n195 = I2[3];
  assign n196 = I2[4];
  assign n197 = I2[5];
  assign n198 = I2[6];
  assign n199 = I2[7];
  assign n200 = I2[8];
  assign n201 = I2[9];
  assign n206 = I1[0];
  assign n207 = I1[1];

  NR2 U82 ( .A(n119), .B(n124), .Z(n73) );
  NR2 U86 ( .A(n125), .B(n132), .Z(n76) );
  NR2 U93 ( .A(n133), .B(n139), .Z(n82) );
  NR2 U111 ( .A(n147), .B(n194), .Z(n98) );
  MUX21L U141 ( .A(n71), .B(n70), .S(n80), .Z(n67) );
  MUX21L U142 ( .A(n73), .B(n74), .S(n77), .Z(n71) );
  MUX21L U143 ( .A(n73), .B(n74), .S(n76), .Z(n70) );
  ND2 U144 ( .A(n119), .B(n124), .Z(n74) );
  ND2 U145 ( .A(n125), .B(n132), .Z(n77) );
  MUX21L U146 ( .A(n209), .B(n210), .S(n80), .Z(O2[4]) );
  EN U147 ( .A(n72), .B(n77), .Z(n209) );
  EN U148 ( .A(n72), .B(n76), .Z(n210) );
  EN U149 ( .A(n119), .B(n124), .Z(n72) );
  FA1A U150 ( .A(n134), .B(n136), .CI(n127), .CO(n124), .S(n125) );
  EN U151 ( .A(n67), .B(n62), .Z(n158) );
  EO U152 ( .A(n118), .B(n113), .Z(n62) );
  OR2 U153 ( .A(n140), .B(n145), .Z(n211) );
  MUX21L U154 ( .A(n82), .B(n83), .S(n84), .Z(n80) );
  ND2 U155 ( .A(n133), .B(n139), .Z(n83) );
  MUX21L U156 ( .A(n212), .B(n211), .S(n213), .Z(n84) );
  FA1A U157 ( .A(n121), .B(n128), .CI(n126), .CO(n118), .S(n119) );
  FA1A U158 ( .A(n137), .B(n135), .CI(n141), .CO(n132), .S(n133) );
  AN2P U159 ( .A(n140), .B(n145), .Z(n212) );
  MUX21L U160 ( .A(n99), .B(n98), .S(n146), .Z(n213) );
  FA1A U161 ( .A(n144), .B(n207), .CI(n142), .CO(n139), .S(n140) );
  FA1A U162 ( .A(n201), .B(n199), .CI(n197), .CO(n128), .S(n129) );
  FA1A U163 ( .A(n131), .B(n195), .CI(n129), .CO(n126), .S(n127) );
  HA1 U164 ( .A(n200), .B(n207), .CO(n130), .S(n131) );
  HA1 U165 ( .A(n198), .B(n201), .CO(n143), .S(n144) );
  FA1A U166 ( .A(n206), .B(n196), .CI(n130), .CO(n122), .S(n123) );
  FA1A U167 ( .A(n196), .B(n194), .CI(n138), .CO(n134), .S(n135) );
  IVDA U168 ( .A(n200), .Y(n138) );
  FA1A U169 ( .A(n199), .B(n197), .CI(n195), .CO(n141), .S(n142) );
  FA1A U170 ( .A(n206), .B(n198), .CI(n143), .CO(n136), .S(n137) );
  FA1A U171 ( .A(n200), .B(n198), .CI(n123), .CO(n120), .S(n121) );
  FA1A U172 ( .A(n200), .B(n196), .CI(n206), .CO(n145), .S(n146) );
  EO3P U173 ( .A(n115), .B(n122), .C(n120), .Z(n113) );
  EO3P U174 ( .A(n199), .B(n197), .C(n117), .Z(n115) );
  EO U175 ( .A(n207), .B(n201), .Z(n117) );
  IVP U176 ( .A(n198), .Z(n147) );
  ND2 U177 ( .A(n147), .B(n194), .Z(n99) );
endmodule


module prime_DW_div_uns_10 ( a, b, quotient, remainder, divide_by_0 );
  input [9:0] a;
  input [1:0] b;
  output [9:0] quotient;
  output [1:0] remainder;
  output divide_by_0;
  wire   \u_div/Adiv3_acc[4] , \u_div/Adiv3_acc[5] , n2, n3, n4, n5, n6;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11;

  prime_add_0_root_add_212_I6_DP_OP_297_0_0 \u_div/add_0_root_add_212_I6_DP_OP_297_0_15  ( 
        .I1(a[9:8]), .I2({a, 1'b0, 1'b0}), .I3(a), .I4(a[9:2]), .I5(a[9:4]), 
        .I6(a[9:6]), .O2({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, \u_div/Adiv3_acc[5] , 
        \u_div/Adiv3_acc[4] , SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11}) );
  EN U1 ( .A(n2), .B(n3), .Z(remainder[1]) );
  IVP U2 ( .A(\u_div/Adiv3_acc[4] ), .Z(n6) );
  EN U3 ( .A(n6), .B(a[0]), .Z(remainder[0]) );
  EO U4 ( .A(n4), .B(a[1]), .Z(n2) );
  EO U5 ( .A(\u_div/Adiv3_acc[5] ), .B(\u_div/Adiv3_acc[4] ), .Z(n3) );
  ND2 U6 ( .A(\u_div/Adiv3_acc[4] ), .B(n5), .Z(n4) );
  IVP U7 ( .A(a[0]), .Z(n5) );
endmodule


module prime ( input_no, clock, reset_n, input_valid, result_ready, is_prime
 );
  input [9:0] input_no;
  input clock, reset_n, input_valid;
  output result_ready, is_prime;
  wire   \state[0] , N0, N1, N35, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N52, n57, n58, n59, n60, \rem_74_2/u_div/BInv[3][13] ,
         \rem_74_2/u_div/BInv[3][12] , \rem_74_2/u_div/BInv[3][11] ,
         \rem_74_2/u_div/BInv[3][10] , \rem_74_2/u_div/BInv[3][9] ,
         \rem_74_2/u_div/BInv[3][8] , \rem_74_2/u_div/BInv[3][7] ,
         \rem_74_2/u_div/BInv[3][6] , \rem_74_2/u_div/BInv[3][5] ,
         \rem_74_2/u_div/BInv[3][4] , \rem_74_2/u_div/BInv[3][3] ,
         \rem_74_2/u_div/BInv[3][2] , \rem_74_2/u_div/BInv[3][1] ,
         \rem_74_2/u_div/BInv[3][0] , \rem_74_2/u_div/BInv[5][14] ,
         \rem_74_2/u_div/BInv[5][13] , \rem_74_2/u_div/BInv[5][12] ,
         \rem_74_2/u_div/BInv[5][11] , \rem_74_2/u_div/BInv[5][10] ,
         \rem_74_2/u_div/BInv[5][9] , \rem_74_2/u_div/BInv[5][8] ,
         \rem_74_2/u_div/BInv[5][7] , \rem_74_2/u_div/BInv[5][6] ,
         \rem_74_2/u_div/BInv[5][5] , \rem_74_2/u_div/BInv[5][4] ,
         \rem_74_2/u_div/BInv[5][3] , \rem_74_2/u_div/BInv[5][2] ,
         \rem_74_2/u_div/BInv[5][1] , \rem_74_2/u_div/BInv[5][0] ,
         \rem_74_2/u_div/BInv[6][14] , \rem_74_2/u_div/BInv[6][13] ,
         \rem_74_2/u_div/BInv[6][12] , \rem_74_2/u_div/BInv[6][11] ,
         \rem_74_2/u_div/BInv[6][10] , \rem_74_2/u_div/BInv[6][9] ,
         \rem_74_2/u_div/BInv[6][8] , \rem_74_2/u_div/BInv[6][7] ,
         \rem_74_2/u_div/BInv[6][6] , \rem_74_2/u_div/BInv[6][5] ,
         \rem_74_2/u_div/BInv[6][4] , \rem_74_2/u_div/BInv[6][3] ,
         \rem_74_2/u_div/BInv[6][2] , \rem_74_2/u_div/BInv[6][1] ,
         \rem_74_2/u_div/BInv[7][14] , \rem_74_2/u_div/BInv[7][13] ,
         \rem_74_2/u_div/BInv[7][12] , \rem_74_2/u_div/BInv[7][11] ,
         \rem_74_2/u_div/BInv[7][10] , \rem_74_2/u_div/BInv[7][9] ,
         \rem_74_2/u_div/BInv[7][8] , \rem_74_2/u_div/BInv[7][7] ,
         \rem_74_2/u_div/BInv[7][6] , \rem_74_2/u_div/BInv[7][5] ,
         \rem_74_2/u_div/BInv[7][4] , \rem_74_2/u_div/BInv[7][3] ,
         \rem_74_2/u_div/BInv[7][2] , \rem_74_2/u_div/BInv[7][1] ,
         \rem_74_2/u_div/BInv[7][0] , \rem_74_2/u_div/PartRem[1][11] ,
         \rem_74_2/u_div/PartRem[1][10] , \rem_74_2/u_div/CryOut[1][3] ,
         \rem_74_2/u_div/CryOut[1][2] , \rem_74_2/u_div/CryOut[1][1] ,
         \rem_74_2/u_div/CryOut[1][0] , \rem_74_2/u_div/CryOut[2][2] ,
         \rem_74_2/u_div/CryOut[2][1] , \rem_74_2/u_div/CryOut[2][0] ,
         \rem_74_2/u_div/CryOut[3][2] , \rem_74_2/u_div/CryOut[3][1] ,
         \rem_74_2/u_div/CryOut[3][0] , \rem_74_2/u_div/CryOut[5][2] ,
         \rem_74_2/u_div/CryOut[5][1] , \rem_74_2/u_div/CryOut[5][0] ,
         \rem_74_2/u_div/CryOut[6][2] , \rem_74_2/u_div/CryOut[6][1] ,
         \rem_74_2/u_div/CryOut[6][0] , \rem_74_2/u_div/CryOut[7][2] ,
         \rem_74_2/u_div/CryOut[7][1] , \rem_74_2/u_div/CryOut[7][0] ,
         \rem_74_2/u_div/SumTmp[1][3][2] , \rem_74_2/u_div/SumTmp[1][3][1] ,
         \rem_74_2/u_div/SumTmp[1][3][0] , \rem_74_2/u_div/SumTmp[1][2][5] ,
         \rem_74_2/u_div/SumTmp[1][2][4] , \rem_74_2/u_div/SumTmp[1][2][3] ,
         \rem_74_2/u_div/SumTmp[1][2][2] , \rem_74_2/u_div/SumTmp[1][2][1] ,
         \rem_74_2/u_div/SumTmp[1][2][0] , \rem_74_2/u_div/SumTmp[1][1][8] ,
         \rem_74_2/u_div/SumTmp[1][1][7] , \rem_74_2/u_div/SumTmp[1][1][6] ,
         \rem_74_2/u_div/SumTmp[1][1][5] , \rem_74_2/u_div/SumTmp[1][1][4] ,
         \rem_74_2/u_div/SumTmp[1][1][3] , \rem_74_2/u_div/SumTmp[1][1][2] ,
         \rem_74_2/u_div/SumTmp[1][1][1] , \rem_74_2/u_div/SumTmp[1][1][0] ,
         \rem_74_2/u_div/SumTmp[1][0][9] , \rem_74_2/u_div/SumTmp[1][0][8] ,
         \rem_74_2/u_div/SumTmp[1][0][7] , \rem_74_2/u_div/SumTmp[1][0][6] ,
         \rem_74_2/u_div/SumTmp[1][0][5] , \rem_74_2/u_div/SumTmp[1][0][4] ,
         \rem_74_2/u_div/SumTmp[1][0][3] , \rem_74_2/u_div/SumTmp[1][0][2] ,
         \rem_74_2/u_div/SumTmp[1][0][1] , \rem_74_2/u_div/SumTmp[1][0][0] ,
         \rem_74_2/u_div/SumTmp[2][2][5] , \rem_74_2/u_div/SumTmp[2][2][4] ,
         \rem_74_2/u_div/SumTmp[2][2][3] , \rem_74_2/u_div/SumTmp[2][2][2] ,
         \rem_74_2/u_div/SumTmp[2][2][1] , \rem_74_2/u_div/SumTmp[2][2][0] ,
         \rem_74_2/u_div/SumTmp[2][1][8] , \rem_74_2/u_div/SumTmp[2][1][7] ,
         \rem_74_2/u_div/SumTmp[2][1][6] , \rem_74_2/u_div/SumTmp[2][1][5] ,
         \rem_74_2/u_div/SumTmp[2][1][4] , \rem_74_2/u_div/SumTmp[2][1][3] ,
         \rem_74_2/u_div/SumTmp[2][1][2] , \rem_74_2/u_div/SumTmp[2][1][1] ,
         \rem_74_2/u_div/SumTmp[2][1][0] , \rem_74_2/u_div/SumTmp[2][0][9] ,
         \rem_74_2/u_div/SumTmp[2][0][8] , \rem_74_2/u_div/SumTmp[2][0][7] ,
         \rem_74_2/u_div/SumTmp[2][0][6] , \rem_74_2/u_div/SumTmp[2][0][5] ,
         \rem_74_2/u_div/SumTmp[2][0][4] , \rem_74_2/u_div/SumTmp[2][0][3] ,
         \rem_74_2/u_div/SumTmp[2][0][2] , \rem_74_2/u_div/SumTmp[2][0][1] ,
         \rem_74_2/u_div/SumTmp[2][0][0] , \rem_74_2/u_div/SumTmp[3][2][5] ,
         \rem_74_2/u_div/SumTmp[3][2][4] , \rem_74_2/u_div/SumTmp[3][2][3] ,
         \rem_74_2/u_div/SumTmp[3][2][2] , \rem_74_2/u_div/SumTmp[3][2][1] ,
         \rem_74_2/u_div/SumTmp[3][2][0] , \rem_74_2/u_div/SumTmp[3][1][8] ,
         \rem_74_2/u_div/SumTmp[3][1][7] , \rem_74_2/u_div/SumTmp[3][1][6] ,
         \rem_74_2/u_div/SumTmp[3][1][5] , \rem_74_2/u_div/SumTmp[3][1][4] ,
         \rem_74_2/u_div/SumTmp[3][1][3] , \rem_74_2/u_div/SumTmp[3][1][2] ,
         \rem_74_2/u_div/SumTmp[3][1][1] , \rem_74_2/u_div/SumTmp[3][1][0] ,
         \rem_74_2/u_div/SumTmp[3][0][9] , \rem_74_2/u_div/SumTmp[3][0][8] ,
         \rem_74_2/u_div/SumTmp[3][0][7] , \rem_74_2/u_div/SumTmp[3][0][6] ,
         \rem_74_2/u_div/SumTmp[3][0][5] , \rem_74_2/u_div/SumTmp[3][0][4] ,
         \rem_74_2/u_div/SumTmp[3][0][3] , \rem_74_2/u_div/SumTmp[3][0][2] ,
         \rem_74_2/u_div/SumTmp[3][0][1] , \rem_74_2/u_div/SumTmp[3][0][0] ,
         \rem_74_2/u_div/SumTmp[4][2][5] , \rem_74_2/u_div/SumTmp[4][2][4] ,
         \rem_74_2/u_div/SumTmp[4][2][3] , \rem_74_2/u_div/SumTmp[4][2][2] ,
         \rem_74_2/u_div/SumTmp[4][2][1] , \rem_74_2/u_div/SumTmp[4][2][0] ,
         \rem_74_2/u_div/SumTmp[4][1][8] , \rem_74_2/u_div/SumTmp[4][1][7] ,
         \rem_74_2/u_div/SumTmp[4][1][6] , \rem_74_2/u_div/SumTmp[4][1][5] ,
         \rem_74_2/u_div/SumTmp[4][1][4] , \rem_74_2/u_div/SumTmp[4][1][3] ,
         \rem_74_2/u_div/SumTmp[4][1][2] , \rem_74_2/u_div/SumTmp[4][1][1] ,
         \rem_74_2/u_div/SumTmp[4][1][0] , \rem_74_2/u_div/SumTmp[4][0][9] ,
         \rem_74_2/u_div/SumTmp[4][0][8] , \rem_74_2/u_div/SumTmp[4][0][7] ,
         \rem_74_2/u_div/SumTmp[4][0][6] , \rem_74_2/u_div/SumTmp[4][0][5] ,
         \rem_74_2/u_div/SumTmp[4][0][4] , \rem_74_2/u_div/SumTmp[4][0][3] ,
         \rem_74_2/u_div/SumTmp[4][0][2] , \rem_74_2/u_div/SumTmp[4][0][1] ,
         \rem_74_2/u_div/SumTmp[4][0][0] , \rem_74_2/u_div/SumTmp[5][2][5] ,
         \rem_74_2/u_div/SumTmp[5][2][4] , \rem_74_2/u_div/SumTmp[5][2][3] ,
         \rem_74_2/u_div/SumTmp[5][2][2] , \rem_74_2/u_div/SumTmp[5][2][1] ,
         \rem_74_2/u_div/SumTmp[5][2][0] , \rem_74_2/u_div/SumTmp[5][1][8] ,
         \rem_74_2/u_div/SumTmp[5][1][7] , \rem_74_2/u_div/SumTmp[5][1][6] ,
         \rem_74_2/u_div/SumTmp[5][1][5] , \rem_74_2/u_div/SumTmp[5][1][4] ,
         \rem_74_2/u_div/SumTmp[5][1][3] , \rem_74_2/u_div/SumTmp[5][1][2] ,
         \rem_74_2/u_div/SumTmp[5][1][1] , \rem_74_2/u_div/SumTmp[5][1][0] ,
         \rem_74_2/u_div/SumTmp[5][0][9] , \rem_74_2/u_div/SumTmp[5][0][8] ,
         \rem_74_2/u_div/SumTmp[5][0][7] , \rem_74_2/u_div/SumTmp[5][0][6] ,
         \rem_74_2/u_div/SumTmp[5][0][5] , \rem_74_2/u_div/SumTmp[5][0][4] ,
         \rem_74_2/u_div/SumTmp[5][0][3] , \rem_74_2/u_div/SumTmp[5][0][2] ,
         \rem_74_2/u_div/SumTmp[5][0][1] , \rem_74_2/u_div/SumTmp[5][0][0] ,
         \rem_74_2/u_div/SumTmp[6][2][5] , \rem_74_2/u_div/SumTmp[6][2][4] ,
         \rem_74_2/u_div/SumTmp[6][2][3] , \rem_74_2/u_div/SumTmp[6][2][2] ,
         \rem_74_2/u_div/SumTmp[6][2][1] , \rem_74_2/u_div/SumTmp[6][2][0] ,
         \rem_74_2/u_div/SumTmp[6][1][8] , \rem_74_2/u_div/SumTmp[6][1][7] ,
         \rem_74_2/u_div/SumTmp[6][1][6] , \rem_74_2/u_div/SumTmp[6][1][5] ,
         \rem_74_2/u_div/SumTmp[6][1][4] , \rem_74_2/u_div/SumTmp[6][1][3] ,
         \rem_74_2/u_div/SumTmp[6][1][2] , \rem_74_2/u_div/SumTmp[6][1][1] ,
         \rem_74_2/u_div/SumTmp[6][1][0] , \rem_74_2/u_div/SumTmp[6][0][9] ,
         \rem_74_2/u_div/SumTmp[6][0][8] , \rem_74_2/u_div/SumTmp[6][0][7] ,
         \rem_74_2/u_div/SumTmp[6][0][6] , \rem_74_2/u_div/SumTmp[6][0][5] ,
         \rem_74_2/u_div/SumTmp[6][0][4] , \rem_74_2/u_div/SumTmp[6][0][3] ,
         \rem_74_2/u_div/SumTmp[6][0][2] , \rem_74_2/u_div/SumTmp[6][0][1] ,
         \rem_74_2/u_div/SumTmp[6][0][0] , \rem_74_2/u_div/SumTmp[7][2][5] ,
         \rem_74_2/u_div/SumTmp[7][2][4] , \rem_74_2/u_div/SumTmp[7][2][3] ,
         \rem_74_2/u_div/SumTmp[7][2][2] , \rem_74_2/u_div/SumTmp[7][2][1] ,
         \rem_74_2/u_div/SumTmp[7][2][0] , \rem_74_2/u_div/SumTmp[7][1][8] ,
         \rem_74_2/u_div/SumTmp[7][1][7] , \rem_74_2/u_div/SumTmp[7][1][6] ,
         \rem_74_2/u_div/SumTmp[7][1][5] , \rem_74_2/u_div/SumTmp[7][1][4] ,
         \rem_74_2/u_div/SumTmp[7][1][3] , \rem_74_2/u_div/SumTmp[7][1][2] ,
         \rem_74_2/u_div/SumTmp[7][1][1] , \rem_74_2/u_div/SumTmp[7][1][0] ,
         \rem_74_2/u_div/SumTmp[7][0][9] , \rem_74_2/u_div/SumTmp[7][0][8] ,
         \rem_74_2/u_div/SumTmp[7][0][7] , \rem_74_2/u_div/SumTmp[7][0][6] ,
         \rem_74_2/u_div/SumTmp[7][0][5] , \rem_74_2/u_div/SumTmp[7][0][4] ,
         \rem_74_2/u_div/SumTmp[7][0][3] , \rem_74_2/u_div/SumTmp[7][0][2] ,
         \rem_74_2/u_div/SumTmp[7][0][1] , \rem_74_2/u_div/SumTmp[7][0][0] ,
         \rem_74_2/quotient[2] , \rem_74_2/quotient[5] ,
         \rem_74_2/quotient[8] , \rem_74/u_div/BInv[3][12] ,
         \rem_74/u_div/BInv[3][11] , \rem_74/u_div/BInv[3][10] ,
         \rem_74/u_div/BInv[3][9] , \rem_74/u_div/BInv[3][8] ,
         \rem_74/u_div/BInv[3][7] , \rem_74/u_div/BInv[3][6] ,
         \rem_74/u_div/BInv[3][5] , \rem_74/u_div/BInv[3][4] ,
         \rem_74/u_div/BInv[3][3] , \rem_74/u_div/BInv[3][2] ,
         \rem_74/u_div/BInv[3][1] , \rem_74/u_div/BInv[3][0] ,
         \rem_74/u_div/BInv[5][13] , \rem_74/u_div/BInv[5][12] ,
         \rem_74/u_div/BInv[5][11] , \rem_74/u_div/BInv[5][10] ,
         \rem_74/u_div/BInv[5][9] , \rem_74/u_div/BInv[5][8] ,
         \rem_74/u_div/BInv[5][7] , \rem_74/u_div/BInv[5][6] ,
         \rem_74/u_div/BInv[5][5] , \rem_74/u_div/BInv[5][4] ,
         \rem_74/u_div/BInv[5][3] , \rem_74/u_div/BInv[5][2] ,
         \rem_74/u_div/BInv[5][1] , \rem_74/u_div/BInv[5][0] ,
         \rem_74/u_div/BInv[6][13] , \rem_74/u_div/BInv[6][12] ,
         \rem_74/u_div/BInv[6][11] , \rem_74/u_div/BInv[6][10] ,
         \rem_74/u_div/BInv[6][9] , \rem_74/u_div/BInv[6][8] ,
         \rem_74/u_div/BInv[6][7] , \rem_74/u_div/BInv[6][6] ,
         \rem_74/u_div/BInv[6][5] , \rem_74/u_div/BInv[6][4] ,
         \rem_74/u_div/BInv[6][3] , \rem_74/u_div/BInv[6][2] ,
         \rem_74/u_div/BInv[6][1] , \rem_74/u_div/BInv[7][13] ,
         \rem_74/u_div/BInv[7][12] , \rem_74/u_div/BInv[7][11] ,
         \rem_74/u_div/BInv[7][10] , \rem_74/u_div/BInv[7][9] ,
         \rem_74/u_div/BInv[7][8] , \rem_74/u_div/BInv[7][7] ,
         \rem_74/u_div/BInv[7][6] , \rem_74/u_div/BInv[7][5] ,
         \rem_74/u_div/BInv[7][4] , \rem_74/u_div/BInv[7][3] ,
         \rem_74/u_div/BInv[7][2] , \rem_74/u_div/BInv[7][1] ,
         \rem_74/u_div/BInv[7][0] , \rem_74/u_div/PartRem[1][11] ,
         \rem_74/u_div/PartRem[1][10] , \rem_74/u_div/CryOut[1][3] ,
         \rem_74/u_div/CryOut[1][2] , \rem_74/u_div/CryOut[1][1] ,
         \rem_74/u_div/CryOut[1][0] , \rem_74/u_div/CryOut[2][2] ,
         \rem_74/u_div/CryOut[2][1] , \rem_74/u_div/CryOut[2][0] ,
         \rem_74/u_div/CryOut[3][2] , \rem_74/u_div/CryOut[3][1] ,
         \rem_74/u_div/CryOut[3][0] , \rem_74/u_div/CryOut[5][2] ,
         \rem_74/u_div/CryOut[5][1] , \rem_74/u_div/CryOut[5][0] ,
         \rem_74/u_div/CryOut[6][2] , \rem_74/u_div/CryOut[6][1] ,
         \rem_74/u_div/CryOut[6][0] , \rem_74/u_div/CryOut[7][2] ,
         \rem_74/u_div/CryOut[7][1] , \rem_74/u_div/CryOut[7][0] ,
         \rem_74/u_div/SumTmp[1][3][2] , \rem_74/u_div/SumTmp[1][3][1] ,
         \rem_74/u_div/SumTmp[1][3][0] , \rem_74/u_div/SumTmp[1][2][5] ,
         \rem_74/u_div/SumTmp[1][2][4] , \rem_74/u_div/SumTmp[1][2][3] ,
         \rem_74/u_div/SumTmp[1][2][2] , \rem_74/u_div/SumTmp[1][2][1] ,
         \rem_74/u_div/SumTmp[1][2][0] , \rem_74/u_div/SumTmp[1][1][8] ,
         \rem_74/u_div/SumTmp[1][1][7] , \rem_74/u_div/SumTmp[1][1][6] ,
         \rem_74/u_div/SumTmp[1][1][5] , \rem_74/u_div/SumTmp[1][1][4] ,
         \rem_74/u_div/SumTmp[1][1][3] , \rem_74/u_div/SumTmp[1][1][2] ,
         \rem_74/u_div/SumTmp[1][1][1] , \rem_74/u_div/SumTmp[1][1][0] ,
         \rem_74/u_div/SumTmp[1][0][9] , \rem_74/u_div/SumTmp[1][0][8] ,
         \rem_74/u_div/SumTmp[1][0][7] , \rem_74/u_div/SumTmp[1][0][6] ,
         \rem_74/u_div/SumTmp[1][0][5] , \rem_74/u_div/SumTmp[1][0][4] ,
         \rem_74/u_div/SumTmp[1][0][3] , \rem_74/u_div/SumTmp[1][0][2] ,
         \rem_74/u_div/SumTmp[1][0][1] , \rem_74/u_div/SumTmp[1][0][0] ,
         \rem_74/u_div/SumTmp[2][2][5] , \rem_74/u_div/SumTmp[2][2][4] ,
         \rem_74/u_div/SumTmp[2][2][3] , \rem_74/u_div/SumTmp[2][2][2] ,
         \rem_74/u_div/SumTmp[2][2][1] , \rem_74/u_div/SumTmp[2][2][0] ,
         \rem_74/u_div/SumTmp[2][1][8] , \rem_74/u_div/SumTmp[2][1][7] ,
         \rem_74/u_div/SumTmp[2][1][6] , \rem_74/u_div/SumTmp[2][1][5] ,
         \rem_74/u_div/SumTmp[2][1][4] , \rem_74/u_div/SumTmp[2][1][3] ,
         \rem_74/u_div/SumTmp[2][1][2] , \rem_74/u_div/SumTmp[2][1][1] ,
         \rem_74/u_div/SumTmp[2][1][0] , \rem_74/u_div/SumTmp[2][0][9] ,
         \rem_74/u_div/SumTmp[2][0][8] , \rem_74/u_div/SumTmp[2][0][7] ,
         \rem_74/u_div/SumTmp[2][0][6] , \rem_74/u_div/SumTmp[2][0][5] ,
         \rem_74/u_div/SumTmp[2][0][4] , \rem_74/u_div/SumTmp[2][0][3] ,
         \rem_74/u_div/SumTmp[2][0][2] , \rem_74/u_div/SumTmp[2][0][1] ,
         \rem_74/u_div/SumTmp[2][0][0] , \rem_74/u_div/SumTmp[3][2][5] ,
         \rem_74/u_div/SumTmp[3][2][4] , \rem_74/u_div/SumTmp[3][2][3] ,
         \rem_74/u_div/SumTmp[3][2][2] , \rem_74/u_div/SumTmp[3][2][1] ,
         \rem_74/u_div/SumTmp[3][2][0] , \rem_74/u_div/SumTmp[3][1][8] ,
         \rem_74/u_div/SumTmp[3][1][7] , \rem_74/u_div/SumTmp[3][1][6] ,
         \rem_74/u_div/SumTmp[3][1][5] , \rem_74/u_div/SumTmp[3][1][4] ,
         \rem_74/u_div/SumTmp[3][1][3] , \rem_74/u_div/SumTmp[3][1][2] ,
         \rem_74/u_div/SumTmp[3][1][1] , \rem_74/u_div/SumTmp[3][1][0] ,
         \rem_74/u_div/SumTmp[3][0][9] , \rem_74/u_div/SumTmp[3][0][8] ,
         \rem_74/u_div/SumTmp[3][0][7] , \rem_74/u_div/SumTmp[3][0][6] ,
         \rem_74/u_div/SumTmp[3][0][5] , \rem_74/u_div/SumTmp[3][0][4] ,
         \rem_74/u_div/SumTmp[3][0][3] , \rem_74/u_div/SumTmp[3][0][2] ,
         \rem_74/u_div/SumTmp[3][0][1] , \rem_74/u_div/SumTmp[3][0][0] ,
         \rem_74/u_div/SumTmp[4][2][5] , \rem_74/u_div/SumTmp[4][2][4] ,
         \rem_74/u_div/SumTmp[4][2][3] , \rem_74/u_div/SumTmp[4][2][2] ,
         \rem_74/u_div/SumTmp[4][2][1] , \rem_74/u_div/SumTmp[4][2][0] ,
         \rem_74/u_div/SumTmp[4][1][8] , \rem_74/u_div/SumTmp[4][1][7] ,
         \rem_74/u_div/SumTmp[4][1][6] , \rem_74/u_div/SumTmp[4][1][5] ,
         \rem_74/u_div/SumTmp[4][1][4] , \rem_74/u_div/SumTmp[4][1][3] ,
         \rem_74/u_div/SumTmp[4][1][2] , \rem_74/u_div/SumTmp[4][1][1] ,
         \rem_74/u_div/SumTmp[4][1][0] , \rem_74/u_div/SumTmp[4][0][9] ,
         \rem_74/u_div/SumTmp[4][0][8] , \rem_74/u_div/SumTmp[4][0][7] ,
         \rem_74/u_div/SumTmp[4][0][6] , \rem_74/u_div/SumTmp[4][0][5] ,
         \rem_74/u_div/SumTmp[4][0][4] , \rem_74/u_div/SumTmp[4][0][3] ,
         \rem_74/u_div/SumTmp[4][0][2] , \rem_74/u_div/SumTmp[4][0][1] ,
         \rem_74/u_div/SumTmp[4][0][0] , \rem_74/u_div/SumTmp[5][2][5] ,
         \rem_74/u_div/SumTmp[5][2][4] , \rem_74/u_div/SumTmp[5][2][3] ,
         \rem_74/u_div/SumTmp[5][2][2] , \rem_74/u_div/SumTmp[5][2][1] ,
         \rem_74/u_div/SumTmp[5][2][0] , \rem_74/u_div/SumTmp[5][1][8] ,
         \rem_74/u_div/SumTmp[5][1][7] , \rem_74/u_div/SumTmp[5][1][6] ,
         \rem_74/u_div/SumTmp[5][1][5] , \rem_74/u_div/SumTmp[5][1][4] ,
         \rem_74/u_div/SumTmp[5][1][3] , \rem_74/u_div/SumTmp[5][1][2] ,
         \rem_74/u_div/SumTmp[5][1][1] , \rem_74/u_div/SumTmp[5][1][0] ,
         \rem_74/u_div/SumTmp[5][0][9] , \rem_74/u_div/SumTmp[5][0][8] ,
         \rem_74/u_div/SumTmp[5][0][7] , \rem_74/u_div/SumTmp[5][0][6] ,
         \rem_74/u_div/SumTmp[5][0][5] , \rem_74/u_div/SumTmp[5][0][4] ,
         \rem_74/u_div/SumTmp[5][0][3] , \rem_74/u_div/SumTmp[5][0][2] ,
         \rem_74/u_div/SumTmp[5][0][1] , \rem_74/u_div/SumTmp[5][0][0] ,
         \rem_74/u_div/SumTmp[6][2][5] , \rem_74/u_div/SumTmp[6][2][4] ,
         \rem_74/u_div/SumTmp[6][2][3] , \rem_74/u_div/SumTmp[6][2][2] ,
         \rem_74/u_div/SumTmp[6][2][1] , \rem_74/u_div/SumTmp[6][2][0] ,
         \rem_74/u_div/SumTmp[6][1][8] , \rem_74/u_div/SumTmp[6][1][7] ,
         \rem_74/u_div/SumTmp[6][1][6] , \rem_74/u_div/SumTmp[6][1][5] ,
         \rem_74/u_div/SumTmp[6][1][4] , \rem_74/u_div/SumTmp[6][1][3] ,
         \rem_74/u_div/SumTmp[6][1][2] , \rem_74/u_div/SumTmp[6][1][1] ,
         \rem_74/u_div/SumTmp[6][1][0] , \rem_74/u_div/SumTmp[6][0][9] ,
         \rem_74/u_div/SumTmp[6][0][8] , \rem_74/u_div/SumTmp[6][0][7] ,
         \rem_74/u_div/SumTmp[6][0][6] , \rem_74/u_div/SumTmp[6][0][5] ,
         \rem_74/u_div/SumTmp[6][0][4] , \rem_74/u_div/SumTmp[6][0][3] ,
         \rem_74/u_div/SumTmp[6][0][2] , \rem_74/u_div/SumTmp[6][0][1] ,
         \rem_74/u_div/SumTmp[6][0][0] , \rem_74/u_div/SumTmp[7][2][5] ,
         \rem_74/u_div/SumTmp[7][2][4] , \rem_74/u_div/SumTmp[7][2][3] ,
         \rem_74/u_div/SumTmp[7][2][2] , \rem_74/u_div/SumTmp[7][2][1] ,
         \rem_74/u_div/SumTmp[7][2][0] , \rem_74/u_div/SumTmp[7][1][8] ,
         \rem_74/u_div/SumTmp[7][1][7] , \rem_74/u_div/SumTmp[7][1][6] ,
         \rem_74/u_div/SumTmp[7][1][5] , \rem_74/u_div/SumTmp[7][1][4] ,
         \rem_74/u_div/SumTmp[7][1][3] , \rem_74/u_div/SumTmp[7][1][2] ,
         \rem_74/u_div/SumTmp[7][1][1] , \rem_74/u_div/SumTmp[7][1][0] ,
         \rem_74/u_div/SumTmp[7][0][9] , \rem_74/u_div/SumTmp[7][0][8] ,
         \rem_74/u_div/SumTmp[7][0][7] , \rem_74/u_div/SumTmp[7][0][6] ,
         \rem_74/u_div/SumTmp[7][0][5] , \rem_74/u_div/SumTmp[7][0][4] ,
         \rem_74/u_div/SumTmp[7][0][3] , \rem_74/u_div/SumTmp[7][0][2] ,
         \rem_74/u_div/SumTmp[7][0][1] , \rem_74/u_div/SumTmp[7][0][0] ,
         \rem_74/quotient[2] , \rem_74/quotient[5] , \rem_74/quotient[8] , n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991;
  wire   [10:0] i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        SYNOPSYS_UNCONNECTED__256, SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, 
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, 
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287, 
        SYNOPSYS_UNCONNECTED__288, SYNOPSYS_UNCONNECTED__289, 
        SYNOPSYS_UNCONNECTED__290, SYNOPSYS_UNCONNECTED__291, 
        SYNOPSYS_UNCONNECTED__292, SYNOPSYS_UNCONNECTED__293, 
        SYNOPSYS_UNCONNECTED__294, SYNOPSYS_UNCONNECTED__295, 
        SYNOPSYS_UNCONNECTED__296, SYNOPSYS_UNCONNECTED__297;

  FD1P \i_reg[10]  ( .D(n983), .CP(clock), .Q(i[10]), .QN(n388) );
  FD1P \i_reg[1]  ( .D(n984), .CP(clock), .Q(i[1]), .QN(n387) );
  FD1P \i_reg[4]  ( .D(n986), .CP(clock), .Q(i[4]), .QN(n375) );
  FD1P \i_reg[5]  ( .D(n987), .CP(clock), .Q(i[5]), .QN(n367) );
  FD1P \i_reg[6]  ( .D(n988), .CP(clock), .Q(i[6]), .QN(n381) );
  FD1P \i_reg[7]  ( .D(n989), .CP(clock), .Q(i[7]), .QN(n385) );
  FD1P \i_reg[8]  ( .D(n990), .CP(clock), .Q(i[8]), .QN(n379) );
  FD1P \i_reg[9]  ( .D(n991), .CP(clock), .Q(i[9]), .QN(n369) );
  prime_DW_mult_uns_0 mult_73 ( .a({n100, n88, n380, n201, n92, n366, n376, 
        n187, n81, n429, n398}), .b({n100, n88, n380, n200, n92, n366, n123, 
        n383, n391, n429, n373}), .product({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, N45, N44, N43, N42, 
        N41, N40, N39, N38, N37, SYNOPSYS_UNCONNECTED__11, N35}) );
  prime_DW01_add_25 \rem_74_2/u_div/u_add_PartRem_2_4  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n975, n974, n394, input_no[8:6]}), 
        .B({1'b1, n198, n115, n168, n413, n400, n401, n420, n270, n417, n409, 
        n429, n178, 1'b1, 1'b1}), .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        \rem_74_2/u_div/SumTmp[4][2][5] , \rem_74_2/u_div/SumTmp[4][2][4] , 
        \rem_74_2/u_div/SumTmp[4][2][3] , \rem_74_2/u_div/SumTmp[4][2][2] , 
        \rem_74_2/u_div/SumTmp[4][2][1] , \rem_74_2/u_div/SumTmp[4][2][0] }), 
        .CO(\rem_74_2/quotient[8] ) );
  prime_DW01_add_74 \rem_74_2/u_div/u_add_PartRem_0_2  ( .A({1'b0, 1'b0, 1'b0, 
        n206, \rem_74_2/u_div/PartRem[1][10] , n960, n959, n957, n955, n954, 
        n953, n952, input_no[2:0]}), .B({1'b1, 1'b1, n300, n267, n112, n76, 
        n197, n401, n420, n290, n417, n409, n429, n178, 1'b1}), .CI(1'b1), 
        .SUM({SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, \rem_74_2/u_div/SumTmp[2][0][9] , 
        \rem_74_2/u_div/SumTmp[2][0][8] , \rem_74_2/u_div/SumTmp[2][0][7] , 
        \rem_74_2/u_div/SumTmp[2][0][6] , \rem_74_2/u_div/SumTmp[2][0][5] , 
        \rem_74_2/u_div/SumTmp[2][0][4] , \rem_74_2/u_div/SumTmp[2][0][3] , 
        \rem_74_2/u_div/SumTmp[2][0][2] , \rem_74_2/u_div/SumTmp[2][0][1] , 
        \rem_74_2/u_div/SumTmp[2][0][0] }), .CO(\rem_74_2/u_div/CryOut[2][0] )
         );
  prime_DW01_add_88 \rem_74_2/u_div/u_add_PartRem_1_7  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, n972, n971, n969, n967, n965, n963, input_no[5:3]}), 
        .B({\rem_74_2/u_div/BInv[7][14] , \rem_74_2/u_div/BInv[7][13] , 
        \rem_74_2/u_div/BInv[7][12] , \rem_74_2/u_div/BInv[7][11] , 
        \rem_74_2/u_div/BInv[7][10] , \rem_74_2/u_div/BInv[7][9] , 
        \rem_74_2/u_div/BInv[7][8] , \rem_74_2/u_div/BInv[7][7] , 
        \rem_74_2/u_div/BInv[7][6] , \rem_74_2/u_div/BInv[7][5] , 
        \rem_74_2/u_div/BInv[7][4] , \rem_74_2/u_div/BInv[7][3] , 
        \rem_74_2/u_div/BInv[7][2] , \rem_74_2/u_div/BInv[7][1] , 
        \rem_74_2/u_div/BInv[7][0] }), .CI(1'b1), .SUM({
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        \rem_74_2/u_div/SumTmp[7][1][8] , \rem_74_2/u_div/SumTmp[7][1][7] , 
        \rem_74_2/u_div/SumTmp[7][1][6] , \rem_74_2/u_div/SumTmp[7][1][5] , 
        \rem_74_2/u_div/SumTmp[7][1][4] , \rem_74_2/u_div/SumTmp[7][1][3] , 
        \rem_74_2/u_div/SumTmp[7][1][2] , \rem_74_2/u_div/SumTmp[7][1][1] , 
        \rem_74_2/u_div/SumTmp[7][1][0] }), .CO(\rem_74_2/u_div/CryOut[7][1] )
         );
  prime_DW01_add_89 \rem_74_2/u_div/u_add_PartRem_1_3  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, n972, n971, n969, n967, n965, n963, input_no[5:3]}), 
        .B({1'b1, \rem_74_2/u_div/BInv[3][13] , \rem_74_2/u_div/BInv[3][12] , 
        \rem_74_2/u_div/BInv[3][11] , \rem_74_2/u_div/BInv[3][10] , 
        \rem_74_2/u_div/BInv[3][9] , \rem_74_2/u_div/BInv[3][8] , 
        \rem_74_2/u_div/BInv[3][7] , \rem_74_2/u_div/BInv[3][6] , 
        \rem_74_2/u_div/BInv[3][5] , \rem_74_2/u_div/BInv[3][4] , 
        \rem_74_2/u_div/BInv[3][3] , \rem_74_2/u_div/BInv[3][2] , 
        \rem_74_2/u_div/BInv[3][1] , \rem_74_2/u_div/BInv[3][0] }), .CI(1'b1), 
        .SUM({SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        \rem_74_2/u_div/SumTmp[3][1][8] , \rem_74_2/u_div/SumTmp[3][1][7] , 
        \rem_74_2/u_div/SumTmp[3][1][6] , \rem_74_2/u_div/SumTmp[3][1][5] , 
        \rem_74_2/u_div/SumTmp[3][1][4] , \rem_74_2/u_div/SumTmp[3][1][3] , 
        \rem_74_2/u_div/SumTmp[3][1][2] , \rem_74_2/u_div/SumTmp[3][1][1] , 
        \rem_74_2/u_div/SumTmp[3][1][0] }), .CO(\rem_74_2/u_div/CryOut[3][1] )
         );
  prime_DW01_add_87 \rem_74_2/u_div/u_add_PartRem_1_5  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, n972, n971, n969, n967, n965, n963, input_no[5:3]}), 
        .B({\rem_74_2/u_div/BInv[5][14] , \rem_74_2/u_div/BInv[5][13] , n188, 
        \rem_74_2/u_div/BInv[5][11] , \rem_74_2/u_div/BInv[5][10] , 
        \rem_74_2/u_div/BInv[5][9] , \rem_74_2/u_div/BInv[5][8] , 
        \rem_74_2/u_div/BInv[5][7] , \rem_74_2/u_div/BInv[5][6] , 
        \rem_74_2/u_div/BInv[5][5] , \rem_74_2/u_div/BInv[5][4] , 
        \rem_74_2/u_div/BInv[5][3] , \rem_74_2/u_div/BInv[5][2] , 
        \rem_74_2/u_div/BInv[5][1] , \rem_74_2/u_div/BInv[5][0] }), .CI(1'b1), 
        .SUM({SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        \rem_74_2/u_div/SumTmp[5][1][8] , \rem_74_2/u_div/SumTmp[5][1][7] , 
        \rem_74_2/u_div/SumTmp[5][1][6] , \rem_74_2/u_div/SumTmp[5][1][5] , 
        \rem_74_2/u_div/SumTmp[5][1][4] , \rem_74_2/u_div/SumTmp[5][1][3] , 
        \rem_74_2/u_div/SumTmp[5][1][2] , \rem_74_2/u_div/SumTmp[5][1][1] , 
        \rem_74_2/u_div/SumTmp[5][1][0] }), .CO(\rem_74_2/u_div/CryOut[5][1] )
         );
  prime_DW01_add_78 \rem_74_2/u_div/u_add_PartRem_1_6  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, n972, n971, n969, n967, n965, n963, input_no[5:3]}), 
        .B({\rem_74_2/u_div/BInv[6][14] , n223, \rem_74_2/u_div/BInv[6][12] , 
        \rem_74_2/u_div/BInv[6][11] , \rem_74_2/u_div/BInv[6][10] , 
        \rem_74_2/u_div/BInv[6][9] , \rem_74_2/u_div/BInv[6][8] , 
        \rem_74_2/u_div/BInv[6][7] , \rem_74_2/u_div/BInv[6][6] , 
        \rem_74_2/u_div/BInv[6][5] , \rem_74_2/u_div/BInv[6][4] , 
        \rem_74_2/u_div/BInv[6][3] , \rem_74_2/u_div/BInv[6][2] , 
        \rem_74_2/u_div/BInv[6][1] , 1'b1}), .CI(1'b1), .SUM({
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        \rem_74_2/u_div/SumTmp[6][1][8] , \rem_74_2/u_div/SumTmp[6][1][7] , 
        \rem_74_2/u_div/SumTmp[6][1][6] , \rem_74_2/u_div/SumTmp[6][1][5] , 
        \rem_74_2/u_div/SumTmp[6][1][4] , \rem_74_2/u_div/SumTmp[6][1][3] , 
        \rem_74_2/u_div/SumTmp[6][1][2] , \rem_74_2/u_div/SumTmp[6][1][1] , 
        \rem_74_2/u_div/SumTmp[6][1][0] }), .CO(\rem_74_2/u_div/CryOut[6][1] )
         );
  prime_DW01_add_76 \rem_74_2/u_div/u_add_PartRem_2_2  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n975, n974, n973, input_no[8:6]}), 
        .B({1'b1, 1'b1, n329, n267, n226, n196, n400, n401, n420, n271, n415, 
        n408, n429, n410, 1'b1}), .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, 
        \rem_74_2/u_div/SumTmp[2][2][5] , \rem_74_2/u_div/SumTmp[2][2][4] , 
        \rem_74_2/u_div/SumTmp[2][2][3] , \rem_74_2/u_div/SumTmp[2][2][2] , 
        \rem_74_2/u_div/SumTmp[2][2][1] , \rem_74_2/u_div/SumTmp[2][2][0] }), 
        .CO(\rem_74_2/u_div/CryOut[2][2] ) );
  prime_DW01_add_97 \rem_74_2/u_div/u_add_PartRem_0_1  ( .A({1'b0, 1'b0, 1'b0, 
        n206, \rem_74_2/u_div/PartRem[1][10] , n960, n958, n957, n955, n954, 
        n953, n952, input_no[2:0]}), .B({1'b1, 1'b1, 1'b1, n198, n267, n168, 
        n196, n197, n146, n420, n290, n417, n409, n429, n176}), .CI(1'b1), 
        .SUM({SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, 
        SYNOPSYS_UNCONNECTED__63, \rem_74_2/u_div/SumTmp[1][0][9] , 
        \rem_74_2/u_div/SumTmp[1][0][8] , \rem_74_2/u_div/SumTmp[1][0][7] , 
        \rem_74_2/u_div/SumTmp[1][0][6] , \rem_74_2/u_div/SumTmp[1][0][5] , 
        \rem_74_2/u_div/SumTmp[1][0][4] , \rem_74_2/u_div/SumTmp[1][0][3] , 
        \rem_74_2/u_div/SumTmp[1][0][2] , \rem_74_2/u_div/SumTmp[1][0][1] , 
        \rem_74_2/u_div/SumTmp[1][0][0] }), .CO(\rem_74_2/u_div/CryOut[1][0] )
         );
  prime_DW01_add_95 \rem_74_2/u_div/u_add_PartRem_0_3  ( .A({1'b0, 1'b0, 1'b0, 
        n206, \rem_74_2/u_div/PartRem[1][10] , n961, n958, n956, n955, n236, 
        n953, n952, input_no[2:0]}), .B({1'b1, \rem_74_2/u_div/BInv[3][13] , 
        \rem_74_2/u_div/BInv[3][12] , \rem_74_2/u_div/BInv[3][11] , n260, 
        \rem_74_2/u_div/BInv[3][9] , \rem_74_2/u_div/BInv[3][8] , 
        \rem_74_2/u_div/BInv[3][7] , \rem_74_2/u_div/BInv[3][6] , 
        \rem_74_2/u_div/BInv[3][5] , \rem_74_2/u_div/BInv[3][4] , 
        \rem_74_2/u_div/BInv[3][3] , \rem_74_2/u_div/BInv[3][2] , 
        \rem_74_2/u_div/BInv[3][1] , \rem_74_2/u_div/BInv[3][0] }), .CI(1'b1), 
        .SUM({SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, \rem_74_2/u_div/SumTmp[3][0][9] , 
        \rem_74_2/u_div/SumTmp[3][0][8] , \rem_74_2/u_div/SumTmp[3][0][7] , 
        \rem_74_2/u_div/SumTmp[3][0][6] , \rem_74_2/u_div/SumTmp[3][0][5] , 
        \rem_74_2/u_div/SumTmp[3][0][4] , \rem_74_2/u_div/SumTmp[3][0][3] , 
        \rem_74_2/u_div/SumTmp[3][0][2] , \rem_74_2/u_div/SumTmp[3][0][1] , 
        \rem_74_2/u_div/SumTmp[3][0][0] }), .CO(\rem_74_2/u_div/CryOut[3][0] )
         );
  prime_DW01_add_98 \rem_74_2/u_div/u_add_PartRem_0_5  ( .A({1'b0, 1'b0, 1'b0, 
        n206, \rem_74_2/u_div/PartRem[1][10] , n960, n958, n957, n955, n236, 
        n953, n952, input_no[2:0]}), .B({\rem_74_2/u_div/BInv[5][14] , 
        \rem_74_2/u_div/BInv[5][13] , n188, \rem_74_2/u_div/BInv[5][11] , 
        \rem_74_2/u_div/BInv[5][10] , \rem_74_2/u_div/BInv[5][9] , 
        \rem_74_2/u_div/BInv[5][8] , \rem_74_2/u_div/BInv[5][7] , 
        \rem_74_2/u_div/BInv[5][6] , \rem_74_2/u_div/BInv[5][5] , 
        \rem_74_2/u_div/BInv[5][4] , \rem_74_2/u_div/BInv[5][3] , 
        \rem_74_2/u_div/BInv[5][2] , \rem_74_2/u_div/BInv[5][1] , 
        \rem_74_2/u_div/BInv[5][0] }), .CI(1'b1), .SUM({
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, 
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        SYNOPSYS_UNCONNECTED__73, \rem_74_2/u_div/SumTmp[5][0][9] , 
        \rem_74_2/u_div/SumTmp[5][0][8] , \rem_74_2/u_div/SumTmp[5][0][7] , 
        \rem_74_2/u_div/SumTmp[5][0][6] , \rem_74_2/u_div/SumTmp[5][0][5] , 
        \rem_74_2/u_div/SumTmp[5][0][4] , \rem_74_2/u_div/SumTmp[5][0][3] , 
        \rem_74_2/u_div/SumTmp[5][0][2] , \rem_74_2/u_div/SumTmp[5][0][1] , 
        \rem_74_2/u_div/SumTmp[5][0][0] }), .CO(\rem_74_2/u_div/CryOut[5][0] )
         );
  prime_DW01_add_82 \rem_74_2/u_div/u_add_PartRem_1_2  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, n972, n971, n969, n967, n965, n963, input_no[5:3]}), 
        .B({1'b1, 1'b1, n300, n267, n112, n76, n400, n401, n420, n270, n415, 
        n408, n429, n176, 1'b1}), .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__74, 
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, 
        SYNOPSYS_UNCONNECTED__79, \rem_74_2/u_div/SumTmp[2][1][8] , 
        \rem_74_2/u_div/SumTmp[2][1][7] , \rem_74_2/u_div/SumTmp[2][1][6] , 
        \rem_74_2/u_div/SumTmp[2][1][5] , \rem_74_2/u_div/SumTmp[2][1][4] , 
        \rem_74_2/u_div/SumTmp[2][1][3] , \rem_74_2/u_div/SumTmp[2][1][2] , 
        \rem_74_2/u_div/SumTmp[2][1][1] , \rem_74_2/u_div/SumTmp[2][1][0] }), 
        .CO(\rem_74_2/u_div/CryOut[2][1] ) );
  prime_DW01_add_79 \rem_74_2/u_div/u_add_PartRem_0_4  ( .A({1'b0, 1'b0, 1'b0, 
        \rem_74_2/u_div/PartRem[1][11] , \rem_74_2/u_div/PartRem[1][10] , n961, 
        n959, n957, n955, n954, n953, n952, input_no[2:0]}), .B({1'b1, n300, 
        n267, n331, n196, n400, n401, n420, n290, n415, n408, n429, n176, 1'b1, 
        1'b1}), .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__80, 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82, 
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        \rem_74_2/u_div/SumTmp[4][0][9] , \rem_74_2/u_div/SumTmp[4][0][8] , 
        \rem_74_2/u_div/SumTmp[4][0][7] , \rem_74_2/u_div/SumTmp[4][0][6] , 
        \rem_74_2/u_div/SumTmp[4][0][5] , \rem_74_2/u_div/SumTmp[4][0][4] , 
        \rem_74_2/u_div/SumTmp[4][0][3] , \rem_74_2/u_div/SumTmp[4][0][2] , 
        \rem_74_2/u_div/SumTmp[4][0][1] , \rem_74_2/u_div/SumTmp[4][0][0] }), 
        .CO(\rem_74_2/quotient[2] ) );
  prime_DW01_add_77 \rem_74_2/u_div/u_add_PartRem_3_1  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        input_no[9]}), .B({1'b1, 1'b1, 1'b1, n329, n933, n226, n232, n979, 
        n980, n159, n270, n416, n976, n427, n410}), .CI(1'b1), .SUM({
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, 
        SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, 
        SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, 
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, 
        SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96, 
        \rem_74_2/u_div/SumTmp[1][3][2] , \rem_74_2/u_div/SumTmp[1][3][1] , 
        \rem_74_2/u_div/SumTmp[1][3][0] }), .CO(\rem_74_2/u_div/CryOut[1][3] )
         );
  prime_DW01_add_56 \rem_74/u_div/u_add_PartRem_2_4  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n949, n948, n947, input_no[8:6]}), .B({
        1'b1, n218, n360, n261, n370, n254, n403, n124, n418, n82, n431, n411, 
        1'b1, 1'b1}), .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, \rem_74/u_div/SumTmp[4][2][5] , 
        \rem_74/u_div/SumTmp[4][2][4] , \rem_74/u_div/SumTmp[4][2][3] , 
        \rem_74/u_div/SumTmp[4][2][2] , \rem_74/u_div/SumTmp[4][2][1] , 
        \rem_74/u_div/SumTmp[4][2][0] }), .CO(\rem_74/quotient[8] ) );
  prime_DW01_add_46 \rem_74/u_div/u_add_PartRem_3_1  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        input_no[9]}), .B({1'b1, 1'b1, 1'b1, n218, n204, n950, n951, n91, n367, 
        n375, n393, n389, n387, n374}), .CI(1'b1), .SUM({
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, 
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, 
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, 
        SYNOPSYS_UNCONNECTED__115, \rem_74/u_div/SumTmp[1][3][2] , 
        \rem_74/u_div/SumTmp[1][3][1] , \rem_74/u_div/SumTmp[1][3][0] }), .CO(
        \rem_74/u_div/CryOut[1][3] ) );
  prime_DW01_add_147 \rem_74/u_div/u_add_PartRem_2_1  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n949, n948, n202, input_no[8:6]}), .B({
        1'b1, 1'b1, 1'b1, n218, n360, n90, n385, n254, n404, n124, n419, n361, 
        n431, n411}), .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, 
        SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, 
        SYNOPSYS_UNCONNECTED__123, \rem_74/u_div/SumTmp[1][2][5] , 
        \rem_74/u_div/SumTmp[1][2][4] , \rem_74/u_div/SumTmp[1][2][3] , 
        \rem_74/u_div/SumTmp[1][2][2] , \rem_74/u_div/SumTmp[1][2][1] , 
        \rem_74/u_div/SumTmp[1][2][0] }), .CO(\rem_74/u_div/CryOut[1][2] ) );
  prime_DW01_add_114 \rem_74/u_div/u_add_PartRem_1_6  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, n946, n945, n944, n942, n214, n174, input_no[5:3]}), .B({
        \rem_74/u_div/BInv[6][13] , \rem_74/u_div/BInv[6][12] , 
        \rem_74/u_div/BInv[6][11] , n245, \rem_74/u_div/BInv[6][9] , 
        \rem_74/u_div/BInv[6][8] , \rem_74/u_div/BInv[6][7] , n243, 
        \rem_74/u_div/BInv[6][5] , \rem_74/u_div/BInv[6][4] , 
        \rem_74/u_div/BInv[6][3] , \rem_74/u_div/BInv[6][2] , 
        \rem_74/u_div/BInv[6][1] , 1'b1}), .CI(1'b1), .SUM({
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, \rem_74/u_div/SumTmp[6][1][8] , 
        \rem_74/u_div/SumTmp[6][1][7] , \rem_74/u_div/SumTmp[6][1][6] , 
        \rem_74/u_div/SumTmp[6][1][5] , \rem_74/u_div/SumTmp[6][1][4] , 
        \rem_74/u_div/SumTmp[6][1][3] , \rem_74/u_div/SumTmp[6][1][2] , 
        \rem_74/u_div/SumTmp[6][1][1] , \rem_74/u_div/SumTmp[6][1][0] }), .CO(
        \rem_74/u_div/CryOut[6][1] ) );
  prime_DW01_add_104 \rem_74/u_div/u_add_PartRem_0_2  ( .A({1'b0, 1'b0, 
        \rem_74/u_div/PartRem[1][11] , \rem_74/u_div/PartRem[1][10] , n941, 
        n940, n316, n938, n937, n936, n935, input_no[2:0]}), .B({1'b1, 1'b1, 
        n101, n89, n90, n370, n254, n404, n405, n419, n82, n430, n178, 1'b1}), 
        .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__129, SYNOPSYS_UNCONNECTED__130, 
        SYNOPSYS_UNCONNECTED__131, SYNOPSYS_UNCONNECTED__132, 
        \rem_74/u_div/SumTmp[2][0][9] , \rem_74/u_div/SumTmp[2][0][8] , 
        \rem_74/u_div/SumTmp[2][0][7] , \rem_74/u_div/SumTmp[2][0][6] , 
        \rem_74/u_div/SumTmp[2][0][5] , \rem_74/u_div/SumTmp[2][0][4] , 
        \rem_74/u_div/SumTmp[2][0][3] , \rem_74/u_div/SumTmp[2][0][2] , 
        \rem_74/u_div/SumTmp[2][0][1] , \rem_74/u_div/SumTmp[2][0][0] }), .CO(
        \rem_74/u_div/CryOut[2][0] ) );
  prime_DW01_add_116 \rem_74/u_div/u_add_PartRem_1_7  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, n946, n333, n944, n291, n211, n174, input_no[5:3]}), .B({
        \rem_74/u_div/BInv[7][13] , \rem_74/u_div/BInv[7][12] , 
        \rem_74/u_div/BInv[7][11] , \rem_74/u_div/BInv[7][10] , n242, 
        \rem_74/u_div/BInv[7][8] , \rem_74/u_div/BInv[7][7] , 
        \rem_74/u_div/BInv[7][6] , n259, \rem_74/u_div/BInv[7][4] , 
        \rem_74/u_div/BInv[7][3] , \rem_74/u_div/BInv[7][2] , 
        \rem_74/u_div/BInv[7][1] , \rem_74/u_div/BInv[7][0] }), .CI(1'b1), 
        .SUM({SYNOPSYS_UNCONNECTED__133, SYNOPSYS_UNCONNECTED__134, 
        SYNOPSYS_UNCONNECTED__135, SYNOPSYS_UNCONNECTED__136, 
        SYNOPSYS_UNCONNECTED__137, \rem_74/u_div/SumTmp[7][1][8] , 
        \rem_74/u_div/SumTmp[7][1][7] , \rem_74/u_div/SumTmp[7][1][6] , 
        \rem_74/u_div/SumTmp[7][1][5] , \rem_74/u_div/SumTmp[7][1][4] , 
        \rem_74/u_div/SumTmp[7][1][3] , \rem_74/u_div/SumTmp[7][1][2] , 
        \rem_74/u_div/SumTmp[7][1][1] , \rem_74/u_div/SumTmp[7][1][0] }), .CO(
        \rem_74/u_div/CryOut[7][1] ) );
  prime_DW01_add_126 \rem_74/u_div/u_add_PartRem_1_5  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, n946, n332, n944, n291, n211, n174, input_no[5:3]}), .B({
        \rem_74/u_div/BInv[5][13] , \rem_74/u_div/BInv[5][12] , 
        \rem_74/u_div/BInv[5][11] , \rem_74/u_div/BInv[5][10] , 
        \rem_74/u_div/BInv[5][9] , \rem_74/u_div/BInv[5][8] , 
        \rem_74/u_div/BInv[5][7] , \rem_74/u_div/BInv[5][6] , 
        \rem_74/u_div/BInv[5][5] , \rem_74/u_div/BInv[5][4] , 
        \rem_74/u_div/BInv[5][3] , \rem_74/u_div/BInv[5][2] , 
        \rem_74/u_div/BInv[5][1] , \rem_74/u_div/BInv[5][0] }), .CI(1'b1), 
        .SUM({SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, \rem_74/u_div/SumTmp[5][1][8] , 
        \rem_74/u_div/SumTmp[5][1][7] , \rem_74/u_div/SumTmp[5][1][6] , 
        \rem_74/u_div/SumTmp[5][1][5] , \rem_74/u_div/SumTmp[5][1][4] , 
        \rem_74/u_div/SumTmp[5][1][3] , \rem_74/u_div/SumTmp[5][1][2] , 
        \rem_74/u_div/SumTmp[5][1][1] , \rem_74/u_div/SumTmp[5][1][0] }), .CO(
        \rem_74/u_div/CryOut[5][1] ) );
  prime_DW01_add_121 \rem_74/u_div/u_add_PartRem_0_7  ( .A({1'b0, 1'b0, 
        \rem_74/u_div/PartRem[1][11] , \rem_74/u_div/PartRem[1][10] , n215, 
        n940, n317, n938, n937, n936, n935, input_no[2:0]}), .B({
        \rem_74/u_div/BInv[7][13] , \rem_74/u_div/BInv[7][12] , 
        \rem_74/u_div/BInv[7][11] , \rem_74/u_div/BInv[7][10] , n251, 
        \rem_74/u_div/BInv[7][8] , \rem_74/u_div/BInv[7][7] , 
        \rem_74/u_div/BInv[7][6] , n259, \rem_74/u_div/BInv[7][4] , 
        \rem_74/u_div/BInv[7][3] , \rem_74/u_div/BInv[7][2] , 
        \rem_74/u_div/BInv[7][1] , \rem_74/u_div/BInv[7][0] }), .CI(1'b1), 
        .SUM({SYNOPSYS_UNCONNECTED__143, SYNOPSYS_UNCONNECTED__144, 
        SYNOPSYS_UNCONNECTED__145, SYNOPSYS_UNCONNECTED__146, 
        \rem_74/u_div/SumTmp[7][0][9] , \rem_74/u_div/SumTmp[7][0][8] , 
        \rem_74/u_div/SumTmp[7][0][7] , \rem_74/u_div/SumTmp[7][0][6] , 
        \rem_74/u_div/SumTmp[7][0][5] , \rem_74/u_div/SumTmp[7][0][4] , 
        \rem_74/u_div/SumTmp[7][0][3] , \rem_74/u_div/SumTmp[7][0][2] , 
        \rem_74/u_div/SumTmp[7][0][1] , \rem_74/u_div/SumTmp[7][0][0] }), .CO(
        \rem_74/u_div/CryOut[7][0] ) );
  prime_DW01_add_123 \rem_74/u_div/u_add_PartRem_0_3  ( .A({1'b0, 1'b0, 
        \rem_74/u_div/PartRem[1][11] , \rem_74/u_div/PartRem[1][10] , n215, 
        n940, n316, n938, n324, n257, n314, input_no[2:0]}), .B({1'b1, 
        \rem_74/u_div/BInv[3][12] , \rem_74/u_div/BInv[3][11] , 
        \rem_74/u_div/BInv[3][10] , n117, \rem_74/u_div/BInv[3][8] , 
        \rem_74/u_div/BInv[3][7] , \rem_74/u_div/BInv[3][6] , n263, n99, 
        \rem_74/u_div/BInv[3][3] , n256, \rem_74/u_div/BInv[3][1] , 
        \rem_74/u_div/BInv[3][0] }), .CI(1'b1), .SUM({
        SYNOPSYS_UNCONNECTED__147, SYNOPSYS_UNCONNECTED__148, 
        SYNOPSYS_UNCONNECTED__149, SYNOPSYS_UNCONNECTED__150, 
        \rem_74/u_div/SumTmp[3][0][9] , \rem_74/u_div/SumTmp[3][0][8] , 
        \rem_74/u_div/SumTmp[3][0][7] , \rem_74/u_div/SumTmp[3][0][6] , 
        \rem_74/u_div/SumTmp[3][0][5] , \rem_74/u_div/SumTmp[3][0][4] , 
        \rem_74/u_div/SumTmp[3][0][3] , \rem_74/u_div/SumTmp[3][0][2] , 
        \rem_74/u_div/SumTmp[3][0][1] , \rem_74/u_div/SumTmp[3][0][0] }), .CO(
        \rem_74/u_div/CryOut[3][0] ) );
  prime_DW01_add_141 \rem_74_2/u_div/u_add_B3  ( .A({1'b1, 1'b1, n329, n115, 
        n226, n413, n362, n401, n159, n271, n417, n408, n429, n411, 1'b1}), 
        .B({1'b1, 1'b1, 1'b1, n330, n148, n331, n413, n400, n401, n420, n271, 
        n415, n409, n427, n386}), .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__151, 
        \rem_74_2/u_div/BInv[3][13] , \rem_74_2/u_div/BInv[3][12] , 
        \rem_74_2/u_div/BInv[3][11] , \rem_74_2/u_div/BInv[3][10] , 
        \rem_74_2/u_div/BInv[3][9] , \rem_74_2/u_div/BInv[3][8] , 
        \rem_74_2/u_div/BInv[3][7] , \rem_74_2/u_div/BInv[3][6] , 
        \rem_74_2/u_div/BInv[3][5] , \rem_74_2/u_div/BInv[3][4] , 
        \rem_74_2/u_div/BInv[3][3] , \rem_74_2/u_div/BInv[3][2] , 
        \rem_74_2/u_div/BInv[3][1] , \rem_74_2/u_div/BInv[3][0] }) );
  prime_DW01_add_111 \rem_74_2/u_div/u_add_PartRem_2_6  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n975, n144, n394, input_no[8:6]}), 
        .B({\rem_74_2/u_div/BInv[6][14] , \rem_74_2/u_div/BInv[6][13] , 
        \rem_74_2/u_div/BInv[6][12] , \rem_74_2/u_div/BInv[6][11] , 
        \rem_74_2/u_div/BInv[6][10] , \rem_74_2/u_div/BInv[6][9] , 
        \rem_74_2/u_div/BInv[6][8] , \rem_74_2/u_div/BInv[6][7] , 
        \rem_74_2/u_div/BInv[6][6] , \rem_74_2/u_div/BInv[6][5] , 
        \rem_74_2/u_div/BInv[6][4] , \rem_74_2/u_div/BInv[6][3] , 
        \rem_74_2/u_div/BInv[6][2] , \rem_74_2/u_div/BInv[6][1] , 1'b1}), .CI(
        1'b1), .SUM({SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, \rem_74_2/u_div/SumTmp[6][2][5] , 
        \rem_74_2/u_div/SumTmp[6][2][4] , \rem_74_2/u_div/SumTmp[6][2][3] , 
        \rem_74_2/u_div/SumTmp[6][2][2] , \rem_74_2/u_div/SumTmp[6][2][1] , 
        \rem_74_2/u_div/SumTmp[6][2][0] }), .CO(\rem_74_2/u_div/CryOut[6][2] )
         );
  prime_DW01_add_138 \rem_74_2/u_div/u_add_PartRem_2_3  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n194, n143, n973, input_no[8:6]}), 
        .B({1'b1, \rem_74_2/u_div/BInv[3][13] , \rem_74_2/u_div/BInv[3][12] , 
        \rem_74_2/u_div/BInv[3][11] , \rem_74_2/u_div/BInv[3][10] , 
        \rem_74_2/u_div/BInv[3][9] , \rem_74_2/u_div/BInv[3][8] , 
        \rem_74_2/u_div/BInv[3][7] , \rem_74_2/u_div/BInv[3][6] , 
        \rem_74_2/u_div/BInv[3][5] , \rem_74_2/u_div/BInv[3][4] , 
        \rem_74_2/u_div/BInv[3][3] , \rem_74_2/u_div/BInv[3][2] , 
        \rem_74_2/u_div/BInv[3][1] , \rem_74_2/u_div/BInv[3][0] }), .CI(1'b1), 
        .SUM({SYNOPSYS_UNCONNECTED__161, SYNOPSYS_UNCONNECTED__162, 
        SYNOPSYS_UNCONNECTED__163, SYNOPSYS_UNCONNECTED__164, 
        SYNOPSYS_UNCONNECTED__165, SYNOPSYS_UNCONNECTED__166, 
        SYNOPSYS_UNCONNECTED__167, SYNOPSYS_UNCONNECTED__168, 
        SYNOPSYS_UNCONNECTED__169, \rem_74_2/u_div/SumTmp[3][2][5] , 
        \rem_74_2/u_div/SumTmp[3][2][4] , \rem_74_2/u_div/SumTmp[3][2][3] , 
        \rem_74_2/u_div/SumTmp[3][2][2] , \rem_74_2/u_div/SumTmp[3][2][1] , 
        \rem_74_2/u_div/SumTmp[3][2][0] }), .CO(\rem_74_2/u_div/CryOut[3][2] )
         );
  prime_DW01_add_100 \rem_74/u_div/u_add_PartRem_0_4  ( .A({1'b0, 1'b0, 
        \rem_74/u_div/PartRem[1][11] , \rem_74/u_div/PartRem[1][10] , n941, 
        n940, n939, n938, n157, n257, n209, input_no[2:0]}), .B({1'b1, n101, 
        n89, n261, n372, n254, n404, n407, n419, n82, n432, n176, 1'b1, 1'b1}), 
        .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        \rem_74/u_div/SumTmp[4][0][9] , \rem_74/u_div/SumTmp[4][0][8] , 
        \rem_74/u_div/SumTmp[4][0][7] , \rem_74/u_div/SumTmp[4][0][6] , 
        \rem_74/u_div/SumTmp[4][0][5] , \rem_74/u_div/SumTmp[4][0][4] , 
        \rem_74/u_div/SumTmp[4][0][3] , \rem_74/u_div/SumTmp[4][0][2] , 
        \rem_74/u_div/SumTmp[4][0][1] , \rem_74/u_div/SumTmp[4][0][0] }), .CO(
        \rem_74/quotient[2] ) );
  prime_DW01_add_149 \rem_74/u_div/u_add_PartRem_2_2  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n949, n948, n203, input_no[8:6]}), .B({
        1'b1, 1'b1, n218, n360, n261, n372, n254, n403, n124, n419, n361, n430, 
        n411, 1'b1}), .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__174, 
        SYNOPSYS_UNCONNECTED__175, SYNOPSYS_UNCONNECTED__176, 
        SYNOPSYS_UNCONNECTED__177, SYNOPSYS_UNCONNECTED__178, 
        SYNOPSYS_UNCONNECTED__179, SYNOPSYS_UNCONNECTED__180, 
        SYNOPSYS_UNCONNECTED__181, \rem_74/u_div/SumTmp[2][2][5] , 
        \rem_74/u_div/SumTmp[2][2][4] , \rem_74/u_div/SumTmp[2][2][3] , 
        \rem_74/u_div/SumTmp[2][2][2] , \rem_74/u_div/SumTmp[2][2][1] , 
        \rem_74/u_div/SumTmp[2][2][0] }), .CO(\rem_74/u_div/CryOut[2][2] ) );
  prime_DW01_add_134 \rem_74/u_div/u_add_PartRem_0_5  ( .A({1'b0, 1'b0, 
        \rem_74/u_div/PartRem[1][11] , \rem_74/u_div/PartRem[1][10] , n215, 
        n239, n317, n938, n324, n165, n126, input_no[2:0]}), .B({
        \rem_74/u_div/BInv[5][13] , \rem_74/u_div/BInv[5][12] , 
        \rem_74/u_div/BInv[5][11] , n127, \rem_74/u_div/BInv[5][9] , 
        \rem_74/u_div/BInv[5][8] , \rem_74/u_div/BInv[5][7] , 
        \rem_74/u_div/BInv[5][6] , \rem_74/u_div/BInv[5][5] , 
        \rem_74/u_div/BInv[5][4] , \rem_74/u_div/BInv[5][3] , 
        \rem_74/u_div/BInv[5][2] , \rem_74/u_div/BInv[5][1] , 
        \rem_74/u_div/BInv[5][0] }), .CI(1'b1), .SUM({
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        \rem_74/u_div/SumTmp[5][0][9] , \rem_74/u_div/SumTmp[5][0][8] , 
        \rem_74/u_div/SumTmp[5][0][7] , \rem_74/u_div/SumTmp[5][0][6] , 
        \rem_74/u_div/SumTmp[5][0][5] , \rem_74/u_div/SumTmp[5][0][4] , 
        \rem_74/u_div/SumTmp[5][0][3] , \rem_74/u_div/SumTmp[5][0][2] , 
        \rem_74/u_div/SumTmp[5][0][1] , \rem_74/u_div/SumTmp[5][0][0] }), .CO(
        \rem_74/u_div/CryOut[5][0] ) );
  prime_DW01_add_133 \rem_74/u_div/u_add_PartRem_0_1  ( .A({1'b0, 1'b0, 
        \rem_74/u_div/PartRem[1][11] , \rem_74/u_div/PartRem[1][10] , n941, 
        n940, n317, n938, n324, n165, n126, input_no[2:0]}), .B({1'b1, 1'b1, 
        1'b1, n101, n89, n90, n370, n254, n404, n405, n418, n82, n430, n176}), 
        .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        \rem_74/u_div/SumTmp[1][0][9] , \rem_74/u_div/SumTmp[1][0][8] , 
        \rem_74/u_div/SumTmp[1][0][7] , \rem_74/u_div/SumTmp[1][0][6] , 
        \rem_74/u_div/SumTmp[1][0][5] , \rem_74/u_div/SumTmp[1][0][4] , 
        \rem_74/u_div/SumTmp[1][0][3] , \rem_74/u_div/SumTmp[1][0][2] , 
        \rem_74/u_div/SumTmp[1][0][1] , \rem_74/u_div/SumTmp[1][0][0] }), .CO(
        \rem_74/u_div/CryOut[1][0] ) );
  prime_DW01_sub_4 \rem_74_2/u_div/u_add_B7  ( .A({n198, n267, n331, n413, 
        n362, n401, n420, n270, n415, n408, n429, n411, 1'b1, 1'b1, 1'b1}), 
        .B({1'b1, 1'b1, 1'b1, n329, n281, n112, n413, n362, n402, n142, n270, 
        n416, n87, n429, n386}), .CI(1'b1), .DIFF({
        \rem_74_2/u_div/BInv[7][14] , \rem_74_2/u_div/BInv[7][13] , 
        \rem_74_2/u_div/BInv[7][12] , \rem_74_2/u_div/BInv[7][11] , 
        \rem_74_2/u_div/BInv[7][10] , \rem_74_2/u_div/BInv[7][9] , 
        \rem_74_2/u_div/BInv[7][8] , \rem_74_2/u_div/BInv[7][7] , 
        \rem_74_2/u_div/BInv[7][6] , \rem_74_2/u_div/BInv[7][5] , 
        \rem_74_2/u_div/BInv[7][4] , \rem_74_2/u_div/BInv[7][3] , 
        \rem_74_2/u_div/BInv[7][2] , \rem_74_2/u_div/BInv[7][1] , 
        \rem_74_2/u_div/BInv[7][0] }) );
  prime_DW01_add_112 \rem_74_2/u_div/u_add_PartRem_0_7  ( .A({1'b0, 1'b0, 1'b0, 
        n206, \rem_74_2/u_div/PartRem[1][10] , n961, n958, n956, n955, n236, 
        n953, n952, input_no[2:0]}), .B({\rem_74_2/u_div/BInv[7][14] , 
        \rem_74_2/u_div/BInv[7][13] , \rem_74_2/u_div/BInv[7][12] , 
        \rem_74_2/u_div/BInv[7][11] , \rem_74_2/u_div/BInv[7][10] , 
        \rem_74_2/u_div/BInv[7][9] , \rem_74_2/u_div/BInv[7][8] , 
        \rem_74_2/u_div/BInv[7][7] , \rem_74_2/u_div/BInv[7][6] , 
        \rem_74_2/u_div/BInv[7][5] , \rem_74_2/u_div/BInv[7][4] , 
        \rem_74_2/u_div/BInv[7][3] , \rem_74_2/u_div/BInv[7][2] , 
        \rem_74_2/u_div/BInv[7][1] , \rem_74_2/u_div/BInv[7][0] }), .CI(1'b1), 
        .SUM({SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, \rem_74_2/u_div/SumTmp[7][0][9] , 
        \rem_74_2/u_div/SumTmp[7][0][8] , \rem_74_2/u_div/SumTmp[7][0][7] , 
        \rem_74_2/u_div/SumTmp[7][0][6] , \rem_74_2/u_div/SumTmp[7][0][5] , 
        \rem_74_2/u_div/SumTmp[7][0][4] , \rem_74_2/u_div/SumTmp[7][0][3] , 
        \rem_74_2/u_div/SumTmp[7][0][2] , \rem_74_2/u_div/SumTmp[7][0][1] , 
        \rem_74_2/u_div/SumTmp[7][0][0] }), .CO(\rem_74_2/u_div/CryOut[7][0] )
         );
  prime_DW01_add_148 \rem_74_2/u_div/u_add_PartRem_2_1  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n975, n143, n973, input_no[8:6]}), 
        .B({1'b1, 1'b1, 1'b1, n198, n267, n168, n76, n362, n401, n420, n270, 
        n417, n409, n429, n386}), .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        \rem_74_2/u_div/SumTmp[1][2][5] , \rem_74_2/u_div/SumTmp[1][2][4] , 
        \rem_74_2/u_div/SumTmp[1][2][3] , \rem_74_2/u_div/SumTmp[1][2][2] , 
        \rem_74_2/u_div/SumTmp[1][2][1] , \rem_74_2/u_div/SumTmp[1][2][0] }), 
        .CO(\rem_74_2/u_div/CryOut[1][2] ) );
  prime_DW01_add_154 \rem_74/u_div/u_add_PartRem_2_3  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n949, n948, n202, input_no[8:6]}), .B({
        1'b1, \rem_74/u_div/BInv[3][12] , \rem_74/u_div/BInv[3][11] , 
        \rem_74/u_div/BInv[3][10] , \rem_74/u_div/BInv[3][9] , 
        \rem_74/u_div/BInv[3][8] , \rem_74/u_div/BInv[3][7] , 
        \rem_74/u_div/BInv[3][6] , \rem_74/u_div/BInv[3][5] , 
        \rem_74/u_div/BInv[3][4] , \rem_74/u_div/BInv[3][3] , 
        \rem_74/u_div/BInv[3][2] , \rem_74/u_div/BInv[3][1] , 
        \rem_74/u_div/BInv[3][0] }), .CI(1'b1), .SUM({
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        \rem_74/u_div/SumTmp[3][2][5] , \rem_74/u_div/SumTmp[3][2][4] , 
        \rem_74/u_div/SumTmp[3][2][3] , \rem_74/u_div/SumTmp[3][2][2] , 
        \rem_74/u_div/SumTmp[3][2][1] , \rem_74/u_div/SumTmp[3][2][0] }), .CO(
        \rem_74/u_div/CryOut[3][2] ) );
  prime_DW01_add_167 \rem_74/u_div/u_add_PartRem_2_5  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n949, n948, n202, input_no[8:6]}), .B({
        \rem_74/u_div/BInv[5][13] , \rem_74/u_div/BInv[5][12] , 
        \rem_74/u_div/BInv[5][11] , \rem_74/u_div/BInv[5][10] , 
        \rem_74/u_div/BInv[5][9] , \rem_74/u_div/BInv[5][8] , 
        \rem_74/u_div/BInv[5][7] , \rem_74/u_div/BInv[5][6] , 
        \rem_74/u_div/BInv[5][5] , \rem_74/u_div/BInv[5][4] , 
        \rem_74/u_div/BInv[5][3] , \rem_74/u_div/BInv[5][2] , 
        \rem_74/u_div/BInv[5][1] , \rem_74/u_div/BInv[5][0] }), .CI(1'b1), 
        .SUM({SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        \rem_74/u_div/SumTmp[5][2][5] , \rem_74/u_div/SumTmp[5][2][4] , 
        \rem_74/u_div/SumTmp[5][2][3] , \rem_74/u_div/SumTmp[5][2][2] , 
        \rem_74/u_div/SumTmp[5][2][1] , \rem_74/u_div/SumTmp[5][2][0] }), .CO(
        \rem_74/u_div/CryOut[5][2] ) );
  prime_DW01_add_157 \rem_74/u_div/u_add_PartRem_2_6  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n949, n948, n202, input_no[8:6]}), .B({
        \rem_74/u_div/BInv[6][13] , \rem_74/u_div/BInv[6][12] , 
        \rem_74/u_div/BInv[6][11] , \rem_74/u_div/BInv[6][10] , 
        \rem_74/u_div/BInv[6][9] , \rem_74/u_div/BInv[6][8] , 
        \rem_74/u_div/BInv[6][7] , \rem_74/u_div/BInv[6][6] , 
        \rem_74/u_div/BInv[6][5] , \rem_74/u_div/BInv[6][4] , 
        \rem_74/u_div/BInv[6][3] , \rem_74/u_div/BInv[6][2] , 
        \rem_74/u_div/BInv[6][1] , 1'b1}), .CI(1'b1), .SUM({
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        \rem_74/u_div/SumTmp[6][2][5] , \rem_74/u_div/SumTmp[6][2][4] , 
        \rem_74/u_div/SumTmp[6][2][3] , \rem_74/u_div/SumTmp[6][2][2] , 
        \rem_74/u_div/SumTmp[6][2][1] , \rem_74/u_div/SumTmp[6][2][0] }), .CO(
        \rem_74/u_div/CryOut[6][2] ) );
  prime_DW01_add_156 \rem_74/u_div/u_add_PartRem_1_4  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, n946, n945, n943, n942, n213, n174, input_no[5:3]}), .B({
        1'b1, n101, n360, n90, n372, n254, n404, n406, n419, n361, n431, n178, 
        1'b1, 1'b1}), .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__228, 
        SYNOPSYS_UNCONNECTED__229, SYNOPSYS_UNCONNECTED__230, 
        SYNOPSYS_UNCONNECTED__231, SYNOPSYS_UNCONNECTED__232, 
        \rem_74/u_div/SumTmp[4][1][8] , \rem_74/u_div/SumTmp[4][1][7] , 
        \rem_74/u_div/SumTmp[4][1][6] , \rem_74/u_div/SumTmp[4][1][5] , 
        \rem_74/u_div/SumTmp[4][1][4] , \rem_74/u_div/SumTmp[4][1][3] , 
        \rem_74/u_div/SumTmp[4][1][2] , \rem_74/u_div/SumTmp[4][1][1] , 
        \rem_74/u_div/SumTmp[4][1][0] }), .CO(\rem_74/quotient[5] ) );
  prime_DW01_add_176 \rem_74_2/u_div/u_add_PartRem_2_7  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n194, n144, n973, input_no[8:6]}), 
        .B({\rem_74_2/u_div/BInv[7][14] , \rem_74_2/u_div/BInv[7][13] , 
        \rem_74_2/u_div/BInv[7][12] , \rem_74_2/u_div/BInv[7][11] , 
        \rem_74_2/u_div/BInv[7][10] , \rem_74_2/u_div/BInv[7][9] , 
        \rem_74_2/u_div/BInv[7][8] , \rem_74_2/u_div/BInv[7][7] , 
        \rem_74_2/u_div/BInv[7][6] , \rem_74_2/u_div/BInv[7][5] , 
        \rem_74_2/u_div/BInv[7][4] , \rem_74_2/u_div/BInv[7][3] , 
        \rem_74_2/u_div/BInv[7][2] , \rem_74_2/u_div/BInv[7][1] , 
        \rem_74_2/u_div/BInv[7][0] }), .CI(1'b1), .SUM({
        SYNOPSYS_UNCONNECTED__233, SYNOPSYS_UNCONNECTED__234, 
        SYNOPSYS_UNCONNECTED__235, SYNOPSYS_UNCONNECTED__236, 
        SYNOPSYS_UNCONNECTED__237, SYNOPSYS_UNCONNECTED__238, 
        SYNOPSYS_UNCONNECTED__239, SYNOPSYS_UNCONNECTED__240, 
        SYNOPSYS_UNCONNECTED__241, \rem_74_2/u_div/SumTmp[7][2][5] , 
        \rem_74_2/u_div/SumTmp[7][2][4] , \rem_74_2/u_div/SumTmp[7][2][3] , 
        \rem_74_2/u_div/SumTmp[7][2][2] , \rem_74_2/u_div/SumTmp[7][2][1] , 
        \rem_74_2/u_div/SumTmp[7][2][0] }), .CO(\rem_74_2/u_div/CryOut[7][2] )
         );
  prime_DW01_add_198 \rem_74/u_div/u_add_PartRem_2_7  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n949, n948, n203, input_no[8:6]}), .B({
        \rem_74/u_div/BInv[7][13] , \rem_74/u_div/BInv[7][12] , 
        \rem_74/u_div/BInv[7][11] , \rem_74/u_div/BInv[7][10] , 
        \rem_74/u_div/BInv[7][9] , \rem_74/u_div/BInv[7][8] , 
        \rem_74/u_div/BInv[7][7] , \rem_74/u_div/BInv[7][6] , 
        \rem_74/u_div/BInv[7][5] , \rem_74/u_div/BInv[7][4] , 
        \rem_74/u_div/BInv[7][3] , \rem_74/u_div/BInv[7][2] , 
        \rem_74/u_div/BInv[7][1] , \rem_74/u_div/BInv[7][0] }), .CI(1'b1), 
        .SUM({SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        \rem_74/u_div/SumTmp[7][2][5] , \rem_74/u_div/SumTmp[7][2][4] , 
        \rem_74/u_div/SumTmp[7][2][3] , \rem_74/u_div/SumTmp[7][2][2] , 
        \rem_74/u_div/SumTmp[7][2][1] , \rem_74/u_div/SumTmp[7][2][0] }), .CO(
        \rem_74/u_div/CryOut[7][2] ) );
  prime_DW01_add_204 \rem_74_2/u_div/u_add_PartRem_1_1  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, n972, n971, n969, n967, n965, n963, input_no[5:3]}), 
        .B({1'b1, 1'b1, 1'b1, n330, n267, n168, n196, n197, n401, n420, n290, 
        n415, n408, n429, n178}), .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__250, 
        SYNOPSYS_UNCONNECTED__251, SYNOPSYS_UNCONNECTED__252, 
        SYNOPSYS_UNCONNECTED__253, SYNOPSYS_UNCONNECTED__254, 
        SYNOPSYS_UNCONNECTED__255, \rem_74_2/u_div/SumTmp[1][1][8] , 
        \rem_74_2/u_div/SumTmp[1][1][7] , \rem_74_2/u_div/SumTmp[1][1][6] , 
        \rem_74_2/u_div/SumTmp[1][1][5] , \rem_74_2/u_div/SumTmp[1][1][4] , 
        \rem_74_2/u_div/SumTmp[1][1][3] , \rem_74_2/u_div/SumTmp[1][1][2] , 
        \rem_74_2/u_div/SumTmp[1][1][1] , \rem_74_2/u_div/SumTmp[1][1][0] }), 
        .CO(\rem_74_2/u_div/CryOut[1][1] ) );
  prime_DW01_add_201 \rem_74/u_div/u_add_PartRem_1_1  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, n946, n333, n944, n291, n211, n174, input_no[5:3]}), .B({
        1'b1, 1'b1, 1'b1, n101, n89, n90, n372, n254, n404, n405, n419, n361, 
        n430, n411}), .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__256, 
        SYNOPSYS_UNCONNECTED__257, SYNOPSYS_UNCONNECTED__258, 
        SYNOPSYS_UNCONNECTED__259, SYNOPSYS_UNCONNECTED__260, 
        \rem_74/u_div/SumTmp[1][1][8] , \rem_74/u_div/SumTmp[1][1][7] , 
        \rem_74/u_div/SumTmp[1][1][6] , \rem_74/u_div/SumTmp[1][1][5] , 
        \rem_74/u_div/SumTmp[1][1][4] , \rem_74/u_div/SumTmp[1][1][3] , 
        \rem_74/u_div/SumTmp[1][1][2] , \rem_74/u_div/SumTmp[1][1][1] , 
        \rem_74/u_div/SumTmp[1][1][0] }), .CO(\rem_74/u_div/CryOut[1][1] ) );
  prime_DW01_add_205 \rem_74/u_div/u_add_PartRem_1_3  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, n946, n332, n216, n208, n210, n174, input_no[5:3]}), .B({
        1'b1, \rem_74/u_div/BInv[3][12] , \rem_74/u_div/BInv[3][11] , 
        \rem_74/u_div/BInv[3][10] , \rem_74/u_div/BInv[3][9] , 
        \rem_74/u_div/BInv[3][8] , \rem_74/u_div/BInv[3][7] , 
        \rem_74/u_div/BInv[3][6] , n263, n99, \rem_74/u_div/BInv[3][3] , n256, 
        \rem_74/u_div/BInv[3][1] , \rem_74/u_div/BInv[3][0] }), .CI(1'b1), 
        .SUM({SYNOPSYS_UNCONNECTED__261, SYNOPSYS_UNCONNECTED__262, 
        SYNOPSYS_UNCONNECTED__263, SYNOPSYS_UNCONNECTED__264, 
        SYNOPSYS_UNCONNECTED__265, \rem_74/u_div/SumTmp[3][1][8] , 
        \rem_74/u_div/SumTmp[3][1][7] , \rem_74/u_div/SumTmp[3][1][6] , 
        \rem_74/u_div/SumTmp[3][1][5] , \rem_74/u_div/SumTmp[3][1][4] , 
        \rem_74/u_div/SumTmp[3][1][3] , \rem_74/u_div/SumTmp[3][1][2] , 
        \rem_74/u_div/SumTmp[3][1][1] , \rem_74/u_div/SumTmp[3][1][0] }), .CO(
        \rem_74/u_div/CryOut[3][1] ) );
  prime_DW01_add_203 \rem_74/u_div/u_add_PartRem_1_2  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, n946, n333, n944, n291, n210, n174, input_no[5:3]}), .B({
        1'b1, 1'b1, n101, n360, n261, n371, n254, n404, n407, n419, n82, n430, 
        n410, 1'b1}), .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__266, 
        SYNOPSYS_UNCONNECTED__267, SYNOPSYS_UNCONNECTED__268, 
        SYNOPSYS_UNCONNECTED__269, SYNOPSYS_UNCONNECTED__270, 
        \rem_74/u_div/SumTmp[2][1][8] , \rem_74/u_div/SumTmp[2][1][7] , 
        \rem_74/u_div/SumTmp[2][1][6] , \rem_74/u_div/SumTmp[2][1][5] , 
        \rem_74/u_div/SumTmp[2][1][4] , \rem_74/u_div/SumTmp[2][1][3] , 
        \rem_74/u_div/SumTmp[2][1][2] , \rem_74/u_div/SumTmp[2][1][1] , 
        \rem_74/u_div/SumTmp[2][1][0] }), .CO(\rem_74/u_div/CryOut[2][1] ) );
  prime_DW01_add_232 \rem_74_2/u_div/u_add_B5  ( .A({1'b1, n330, n267, n412, 
        n76, n362, n146, n142, n271, n415, n409, n429, n411, 1'b1, 1'b1}), .B(
        {1'b1, 1'b1, 1'b1, n198, n281, n168, n413, n979, n146, n142, n270, 
        n417, n408, n429, n386}), .CI(1'b1), .SUM({
        \rem_74_2/u_div/BInv[5][14] , \rem_74_2/u_div/BInv[5][13] , 
        \rem_74_2/u_div/BInv[5][12] , \rem_74_2/u_div/BInv[5][11] , 
        \rem_74_2/u_div/BInv[5][10] , \rem_74_2/u_div/BInv[5][9] , 
        \rem_74_2/u_div/BInv[5][8] , \rem_74_2/u_div/BInv[5][7] , 
        \rem_74_2/u_div/BInv[5][6] , \rem_74_2/u_div/BInv[5][5] , 
        \rem_74_2/u_div/BInv[5][4] , \rem_74_2/u_div/BInv[5][3] , 
        \rem_74_2/u_div/BInv[5][2] , \rem_74_2/u_div/BInv[5][1] , 
        \rem_74_2/u_div/BInv[5][0] }) );
  prime_DW01_add_231 \rem_74_2/u_div/u_add_PartRem_2_5  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n194, n144, n973, input_no[8:6]}), 
        .B({\rem_74_2/u_div/BInv[5][14] , \rem_74_2/u_div/BInv[5][13] , 
        \rem_74_2/u_div/BInv[5][12] , \rem_74_2/u_div/BInv[5][11] , 
        \rem_74_2/u_div/BInv[5][10] , \rem_74_2/u_div/BInv[5][9] , 
        \rem_74_2/u_div/BInv[5][8] , \rem_74_2/u_div/BInv[5][7] , 
        \rem_74_2/u_div/BInv[5][6] , \rem_74_2/u_div/BInv[5][5] , 
        \rem_74_2/u_div/BInv[5][4] , \rem_74_2/u_div/BInv[5][3] , 
        \rem_74_2/u_div/BInv[5][2] , \rem_74_2/u_div/BInv[5][1] , 
        \rem_74_2/u_div/BInv[5][0] }), .CI(1'b1), .SUM({
        SYNOPSYS_UNCONNECTED__271, SYNOPSYS_UNCONNECTED__272, 
        SYNOPSYS_UNCONNECTED__273, SYNOPSYS_UNCONNECTED__274, 
        SYNOPSYS_UNCONNECTED__275, SYNOPSYS_UNCONNECTED__276, 
        SYNOPSYS_UNCONNECTED__277, SYNOPSYS_UNCONNECTED__278, 
        SYNOPSYS_UNCONNECTED__279, \rem_74_2/u_div/SumTmp[5][2][5] , 
        \rem_74_2/u_div/SumTmp[5][2][4] , \rem_74_2/u_div/SumTmp[5][2][3] , 
        \rem_74_2/u_div/SumTmp[5][2][2] , \rem_74_2/u_div/SumTmp[5][2][1] , 
        \rem_74_2/u_div/SumTmp[5][2][0] }), .CO(\rem_74_2/u_div/CryOut[5][2] )
         );
  prime_DW01_add_224 \rem_74/u_div/u_add_PartRem_0_6  ( .A({1'b0, 1'b0, 
        \rem_74/u_div/PartRem[1][11] , \rem_74/u_div/PartRem[1][10] , n941, 
        n940, n316, n938, n937, n165, n935, input_no[2:0]}), .B({
        \rem_74/u_div/BInv[6][13] , \rem_74/u_div/BInv[6][12] , n125, n262, 
        \rem_74/u_div/BInv[6][9] , \rem_74/u_div/BInv[6][8] , 
        \rem_74/u_div/BInv[6][7] , n243, \rem_74/u_div/BInv[6][5] , 
        \rem_74/u_div/BInv[6][4] , \rem_74/u_div/BInv[6][3] , 
        \rem_74/u_div/BInv[6][2] , \rem_74/u_div/BInv[6][1] , 1'b1}), .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        \rem_74/u_div/SumTmp[6][0][9] , \rem_74/u_div/SumTmp[6][0][8] , 
        \rem_74/u_div/SumTmp[6][0][7] , \rem_74/u_div/SumTmp[6][0][6] , 
        \rem_74/u_div/SumTmp[6][0][5] , \rem_74/u_div/SumTmp[6][0][4] , 
        \rem_74/u_div/SumTmp[6][0][3] , \rem_74/u_div/SumTmp[6][0][2] , 
        \rem_74/u_div/SumTmp[6][0][1] , \rem_74/u_div/SumTmp[6][0][0] }), .CO(
        \rem_74/u_div/CryOut[6][0] ) );
  prime_DW01_add_223 \rem_74_2/u_div/u_add_PartRem_1_4  ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, n972, n970, n968, n966, n964, n962, input_no[5:3]}), 
        .B({1'b1, n329, n267, n355, n413, n400, n401, n420, n271, n417, n408, 
        n429, n176, 1'b1, 1'b1}), .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__284, 
        SYNOPSYS_UNCONNECTED__285, SYNOPSYS_UNCONNECTED__286, 
        SYNOPSYS_UNCONNECTED__287, SYNOPSYS_UNCONNECTED__288, 
        SYNOPSYS_UNCONNECTED__289, \rem_74_2/u_div/SumTmp[4][1][8] , 
        \rem_74_2/u_div/SumTmp[4][1][7] , \rem_74_2/u_div/SumTmp[4][1][6] , 
        \rem_74_2/u_div/SumTmp[4][1][5] , \rem_74_2/u_div/SumTmp[4][1][4] , 
        \rem_74_2/u_div/SumTmp[4][1][3] , \rem_74_2/u_div/SumTmp[4][1][2] , 
        \rem_74_2/u_div/SumTmp[4][1][1] , \rem_74_2/u_div/SumTmp[4][1][0] }), 
        .CO(\rem_74_2/quotient[5] ) );
  prime_DW01_add_229 \rem_74_2/u_div/u_add_B6  ( .A({1'b1, n330, n281, n226, 
        n413, n362, n402, n160, n271, n416, n408, n427, n411, 1'b1, 1'b1}), 
        .B({1'b1, 1'b1, n330, n977, n412, n414, n362, n980, n160, n269, n416, 
        n976, n427, n411, 1'b1}), .CI(1'b1), .SUM({
        \rem_74_2/u_div/BInv[6][14] , \rem_74_2/u_div/BInv[6][13] , 
        \rem_74_2/u_div/BInv[6][12] , \rem_74_2/u_div/BInv[6][11] , 
        \rem_74_2/u_div/BInv[6][10] , \rem_74_2/u_div/BInv[6][9] , 
        \rem_74_2/u_div/BInv[6][8] , \rem_74_2/u_div/BInv[6][7] , 
        \rem_74_2/u_div/BInv[6][6] , \rem_74_2/u_div/BInv[6][5] , 
        \rem_74_2/u_div/BInv[6][4] , \rem_74_2/u_div/BInv[6][3] , 
        \rem_74_2/u_div/BInv[6][2] , \rem_74_2/u_div/BInv[6][1] , 
        SYNOPSYS_UNCONNECTED__290}) );
  prime_DW01_add_219 \rem_74_2/u_div/u_add_PartRem_0_6  ( .A({1'b0, 1'b0, 1'b0, 
        \rem_74_2/u_div/PartRem[1][11] , \rem_74_2/u_div/PartRem[1][10] , n960, 
        n958, n956, n955, n236, n953, n952, input_no[2:0]}), .B({
        \rem_74_2/u_div/BInv[6][14] , n223, \rem_74_2/u_div/BInv[6][12] , 
        \rem_74_2/u_div/BInv[6][11] , \rem_74_2/u_div/BInv[6][10] , 
        \rem_74_2/u_div/BInv[6][9] , \rem_74_2/u_div/BInv[6][8] , 
        \rem_74_2/u_div/BInv[6][7] , \rem_74_2/u_div/BInv[6][6] , 
        \rem_74_2/u_div/BInv[6][5] , \rem_74_2/u_div/BInv[6][4] , 
        \rem_74_2/u_div/BInv[6][3] , \rem_74_2/u_div/BInv[6][2] , 
        \rem_74_2/u_div/BInv[6][1] , 1'b1}), .CI(1'b1), .SUM({
        SYNOPSYS_UNCONNECTED__291, SYNOPSYS_UNCONNECTED__292, 
        SYNOPSYS_UNCONNECTED__293, SYNOPSYS_UNCONNECTED__294, 
        SYNOPSYS_UNCONNECTED__295, \rem_74_2/u_div/SumTmp[6][0][9] , 
        \rem_74_2/u_div/SumTmp[6][0][8] , \rem_74_2/u_div/SumTmp[6][0][7] , 
        \rem_74_2/u_div/SumTmp[6][0][6] , \rem_74_2/u_div/SumTmp[6][0][5] , 
        \rem_74_2/u_div/SumTmp[6][0][4] , \rem_74_2/u_div/SumTmp[6][0][3] , 
        \rem_74_2/u_div/SumTmp[6][0][2] , \rem_74_2/u_div/SumTmp[6][0][1] , 
        \rem_74_2/u_div/SumTmp[6][0][0] }), .CO(\rem_74_2/u_div/CryOut[6][0] )
         );
  prime_DW01_sub_8 \rem_74/u_div/u_add_B7  ( .A({n218, n360, n90, n371, n255, 
        n80, n170, n186, n392, n432, n411, 1'b1, 1'b1, 1'b1}), .B({1'b1, 1'b1, 
        1'b1, n218, n369, n379, n371, n381, n367, n93, n393, n390, n428, n397}), .CI(1'b1), .DIFF({\rem_74/u_div/BInv[7][13] , \rem_74/u_div/BInv[7][12] , 
        \rem_74/u_div/BInv[7][11] , \rem_74/u_div/BInv[7][10] , 
        \rem_74/u_div/BInv[7][9] , \rem_74/u_div/BInv[7][8] , 
        \rem_74/u_div/BInv[7][7] , \rem_74/u_div/BInv[7][6] , 
        \rem_74/u_div/BInv[7][5] , \rem_74/u_div/BInv[7][4] , 
        \rem_74/u_div/BInv[7][3] , \rem_74/u_div/BInv[7][2] , 
        \rem_74/u_div/BInv[7][1] , \rem_74/u_div/BInv[7][0] }) );
  prime_DW01_add_240 \rem_74/u_div/u_add_B5  ( .A({1'b1, n101, n360, n90, n371, 
        n381, n80, n351, n113, n390, n85, n397, 1'b1, 1'b1}), .B({1'b1, 1'b1, 
        1'b1, n218, n369, n90, n385, n255, n80, n351, n113, n390, n432, n411}), 
        .CI(1'b1), .SUM({\rem_74/u_div/BInv[5][13] , 
        \rem_74/u_div/BInv[5][12] , \rem_74/u_div/BInv[5][11] , 
        \rem_74/u_div/BInv[5][10] , \rem_74/u_div/BInv[5][9] , 
        \rem_74/u_div/BInv[5][8] , \rem_74/u_div/BInv[5][7] , 
        \rem_74/u_div/BInv[5][6] , \rem_74/u_div/BInv[5][5] , 
        \rem_74/u_div/BInv[5][4] , \rem_74/u_div/BInv[5][3] , 
        \rem_74/u_div/BInv[5][2] , \rem_74/u_div/BInv[5][1] , 
        \rem_74/u_div/BInv[5][0] }) );
  prime_DW01_add_215 \rem_74/u_div/u_add_B6  ( .A({1'b1, n101, n360, n90, n370, 
        n91, n80, n93, n384, n181, n192, n397, 1'b1, 1'b1}), .B({1'b1, 1'b1, 
        n218, n360, n379, n385, n91, n80, n375, n384, n390, n192, n386, 1'b1}), 
        .CI(1'b1), .SUM({\rem_74/u_div/BInv[6][13] , 
        \rem_74/u_div/BInv[6][12] , \rem_74/u_div/BInv[6][11] , 
        \rem_74/u_div/BInv[6][10] , \rem_74/u_div/BInv[6][9] , 
        \rem_74/u_div/BInv[6][8] , \rem_74/u_div/BInv[6][7] , 
        \rem_74/u_div/BInv[6][6] , \rem_74/u_div/BInv[6][5] , 
        \rem_74/u_div/BInv[6][4] , \rem_74/u_div/BInv[6][3] , 
        \rem_74/u_div/BInv[6][2] , \rem_74/u_div/BInv[6][1] , 
        SYNOPSYS_UNCONNECTED__296}) );
  prime_DW01_add_217 \rem_74/u_div/u_add_B3  ( .A({1'b1, 1'b1, n101, n360, 
        n261, n372, n91, n367, n421, n384, n181, n85, n397, 1'b1}), .B({1'b1, 
        1'b1, 1'b1, n218, n360, n90, n385, n381, n80, n421, n384, n389, n192, 
        n411}), .CI(1'b1), .SUM({SYNOPSYS_UNCONNECTED__297, 
        \rem_74/u_div/BInv[3][12] , \rem_74/u_div/BInv[3][11] , 
        \rem_74/u_div/BInv[3][10] , \rem_74/u_div/BInv[3][9] , 
        \rem_74/u_div/BInv[3][8] , \rem_74/u_div/BInv[3][7] , 
        \rem_74/u_div/BInv[3][6] , \rem_74/u_div/BInv[3][5] , 
        \rem_74/u_div/BInv[3][4] , \rem_74/u_div/BInv[3][3] , 
        \rem_74/u_div/BInv[3][2] , \rem_74/u_div/BInv[3][1] , 
        \rem_74/u_div/BInv[3][0] }) );
  FD1P \i_reg[0]  ( .D(n60), .CP(clock), .Q(N52), .QN(n397) );
  FD1P \i_reg[2]  ( .D(n59), .CP(clock), .Q(i[2]), .QN(n390) );
  prime_DW_div_uns_10 rem_65_2 ( .a(input_no), .b({1'b1, 1'b1}), .remainder({
        N1, N0}) );
  FD2 is_prime_reg ( .D(n58), .CP(clock), .CD(reset_n), .Q(is_prime) );
  FD2 result_ready_reg ( .D(n57), .CP(clock), .CD(reset_n), .Q(result_ready), 
        .QN(n931) );
  FD1P \i_reg[3]  ( .D(n985), .CP(clock), .Q(i[3]), .QN(n393) );
  FD2 \state_reg[0]  ( .D(n934), .CP(clock), .CD(reset_n), .Q(\state[0] ), 
        .QN(n932) );
  OR2 U62 ( .A(n312), .B(\rem_74/u_div/CryOut[6][0] ), .Z(n150) );
  IVAP U63 ( .A(n828), .Z(n827) );
  IVP U64 ( .A(n149), .Z(n154) );
  IV U65 ( .A(\rem_74_2/u_div/SumTmp[2][0][8] ), .Z(n191) );
  NR3P U66 ( .A(n199), .B(n284), .C(n498), .Z(n62) );
  B3IP U67 ( .A(n166), .Z2(n416) );
  IVAP U68 ( .A(\rem_74_2/quotient[2] ), .Z(n119) );
  B4I U69 ( .A(n638), .Z(n949) );
  B3I U70 ( .A(n121), .Z1(n115) );
  B4I U71 ( .A(n75), .Z(n196) );
  B3IP U72 ( .A(n240), .Z1(n63), .Z2(n64) );
  B4I U73 ( .A(n690), .Z(n174) );
  B2I U74 ( .A(\rem_74/quotient[5] ), .Z1(n65), .Z2(n66) );
  B5I U75 ( .A(n322), .Z(n215) );
  IVDA U76 ( .A(n298), .Y(n67), .Z(n68) );
  B5I U77 ( .A(n773), .Z(n152) );
  IVDAP U78 ( .A(\rem_74/u_div/CryOut[6][0] ), .Y(n69), .Z(n70) );
  AN2P U79 ( .A(n593), .B(n592), .Z(n71) );
  B3I U80 ( .A(n119), .Z1(n72), .Z2(n73) );
  B3IP U81 ( .A(n87), .Z2(n408) );
  IVDAP U82 ( .A(\rem_74/u_div/CryOut[6][1] ), .Y(n283), .Z(n294) );
  IVP U83 ( .A(\rem_74/u_div/CryOut[6][1] ), .Z(n699) );
  AN3P U84 ( .A(\rem_74/u_div/CryOut[7][1] ), .B(\rem_74/u_div/CryOut[6][1] ), 
        .C(\rem_74/quotient[5] ), .Z(n704) );
  AN2 U85 ( .A(\rem_74_2/u_div/SumTmp[4][1][0] ), .B(n297), .Z(n219) );
  IVP U86 ( .A(n241), .Z(n175) );
  IV U87 ( .A(n427), .Z(n431) );
  B5I U88 ( .A(n319), .Z(n297) );
  B3I U89 ( .A(n93), .Z1(n123), .Z2(n170) );
  IVAP U90 ( .A(n123), .Z(n124) );
  B5I U91 ( .A(n94), .Z(n421) );
  B2I U92 ( .A(n170), .Z1(n377), .Z2(n406) );
  B2I U93 ( .A(n170), .Z1(n376), .Z2(n407) );
  B2I U94 ( .A(n170), .Z1(n378), .Z2(n405) );
  AO2 U95 ( .A(\rem_74/u_div/SumTmp[5][2][3] ), .B(n64), .C(
        \rem_74/u_div/SumTmp[1][2][3] ), .D(n280), .Z(n658) );
  B3I U96 ( .A(\rem_74/u_div/CryOut[2][1] ), .Z1(n235), .Z2(n282) );
  IVA U97 ( .A(n702), .Z(n141) );
  NR3P U98 ( .A(n704), .B(n703), .C(n702), .Z(n74) );
  B5I U99 ( .A(n75), .Z(n76) );
  OR2 U100 ( .A(n679), .B(n678), .Z(n299) );
  MUX21L U101 ( .A(n278), .B(n279), .S(n424), .Z(n579) );
  IVAP U102 ( .A(input_no[9]), .Z(n252) );
  IVA U103 ( .A(\rem_74_2/u_div/CryOut[7][1] ), .Z(n279) );
  B5IP U104 ( .A(i[10]), .Z(n218) );
  IVP U105 ( .A(n195), .Z(n269) );
  AO2 U106 ( .A(\rem_74_2/u_div/SumTmp[4][1][6] ), .B(n338), .C(n128), .D(n246), .Z(n593) );
  AO6 U107 ( .A(\rem_74_2/u_div/SumTmp[4][1][3] ), .B(n338), .C(n611), .Z(n614) );
  IVDA U108 ( .A(n362), .Z(n197) );
  ND2 U109 ( .A(n873), .B(n872), .Z(n877) );
  ND2 U110 ( .A(n879), .B(n878), .Z(n883) );
  IVP U111 ( .A(n81), .Z(n361) );
  IVA U112 ( .A(n920), .Z(n833) );
  IVP U113 ( .A(\rem_74/u_div/SumTmp[7][0][2] ), .Z(n275) );
  IVP U114 ( .A(\rem_74/u_div/SumTmp[3][0][2] ), .Z(n274) );
  IVA U115 ( .A(\rem_74/u_div/SumTmp[7][0][3] ), .Z(n277) );
  IVA U116 ( .A(\rem_74/u_div/SumTmp[3][0][3] ), .Z(n276) );
  IVP U117 ( .A(input_valid), .Z(n289) );
  B4I U118 ( .A(N52), .Z(n374) );
  B3IP U119 ( .A(\rem_74_2/quotient[8] ), .Z1(n78), .Z2(n79) );
  IVP U120 ( .A(n379), .Z(n380) );
  B3I U121 ( .A(n111), .Z1(n81), .Z2(n82) );
  B2I U122 ( .A(n951), .Z1(n200), .Z2(n370) );
  IVDAP U123 ( .A(n387), .Y(n84), .Z(n85) );
  AN2 U124 ( .A(\rem_74_2/quotient[2] ), .B(n110), .Z(n86) );
  ENP U125 ( .A(i[2]), .B(i[1]), .Z(n87) );
  B3IP U126 ( .A(i[5]), .Z1(n80), .Z2(n77) );
  IVA U127 ( .A(\rem_74/u_div/SumTmp[1][3][0] ), .Z(n98) );
  IVP U128 ( .A(input_no[6]), .Z(n434) );
  IVP U129 ( .A(input_no[3]), .Z(n433) );
  IVDA U130 ( .A(n360), .Y(n88), .Z(n89) );
  B4I U131 ( .A(n660), .Z(n944) );
  B3IP U132 ( .A(n950), .Z2(n90) );
  B3IP U133 ( .A(i[6]), .Z1(n91), .Z2(n92) );
  IVDAP U134 ( .A(i[4]), .Y(n93), .Z(n94) );
  AN2P U135 ( .A(n334), .B(n363), .Z(n95) );
  AN2P U136 ( .A(n119), .B(n899), .Z(n96) );
  ND3 U137 ( .A(\rem_74/u_div/CryOut[1][1] ), .B(n235), .C(n158), .Z(n97) );
  IVP U138 ( .A(input_no[8]), .Z(n436) );
  IVDAP U139 ( .A(\rem_74/u_div/BInv[3][4] ), .Z(n99) );
  IVDAP U140 ( .A(n388), .Y(n100), .Z(n101) );
  AN2P U141 ( .A(n464), .B(n912), .Z(n102) );
  IVAP U142 ( .A(n544), .Z(n566) );
  IVAP U143 ( .A(n426), .Z(n103) );
  IVAP U144 ( .A(n426), .Z(n425) );
  IVA U145 ( .A(n308), .Z(n104) );
  IVDA U146 ( .A(n628), .Z(n105) );
  IV U147 ( .A(n899), .Z(n106) );
  B4I U148 ( .A(n581), .Z(n107) );
  IVP U149 ( .A(n581), .Z(n637) );
  AN2P U150 ( .A(n591), .B(n590), .Z(n108) );
  IVDAP U151 ( .A(\rem_74_2/u_div/CryOut[6][0] ), .Y(n110), .Z(n109) );
  IV U152 ( .A(n391), .Z(n111) );
  IVAP U153 ( .A(n167), .Z(n112) );
  IVA U154 ( .A(i[3]), .Z(n113) );
  ND2 U155 ( .A(i[3]), .B(i[2]), .Z(n114) );
  ND2 U156 ( .A(i[3]), .B(i[2]), .Z(n499) );
  B5IP U157 ( .A(n427), .Z(n432) );
  AO2 U158 ( .A(\rem_74/u_div/SumTmp[4][2][3] ), .B(n64), .C(n203), .D(n280), 
        .Z(n654) );
  B3IP U159 ( .A(n355), .Z1(n167), .Z2(n412) );
  IVAP U160 ( .A(n63), .Z(n265) );
  IVP U161 ( .A(n313), .Z(n314) );
  IVDAP U162 ( .A(n241), .Y(n221), .Z(n328) );
  IVDAP U163 ( .A(n771), .Y(n935), .Z(n313) );
  B4I U164 ( .A(n504), .Z(n975) );
  OR2P U165 ( .A(n508), .B(n264), .Z(n506) );
  IVAP U166 ( .A(n559), .Z(n568) );
  IVAP U167 ( .A(n555), .Z(n569) );
  B2I U168 ( .A(n384), .Z1(n187), .Z2(n186) );
  IVA U169 ( .A(n258), .Z(n195) );
  ND4P U170 ( .A(n500), .B(i[7]), .C(i[6]), .D(i[8]), .Z(n498) );
  AN2 U171 ( .A(n334), .B(n655), .Z(n116) );
  IVDA U172 ( .A(\rem_74/u_div/BInv[3][9] ), .Z(n117) );
  AN2P U173 ( .A(n518), .B(n78), .Z(n304) );
  ND2 U174 ( .A(n334), .B(n655), .Z(n118) );
  IVP U175 ( .A(n391), .Z(n392) );
  AO7P U176 ( .A(n855), .B(n854), .C(n853), .Z(n890) );
  IV U177 ( .A(n369), .Z(n120) );
  IV U178 ( .A(n682), .Z(n684) );
  B2I U179 ( .A(n80), .Z1(n366), .Z2(n403) );
  MUX21LP U180 ( .A(n640), .B(n98), .S(\rem_74/u_div/CryOut[1][3] ), .Z(n947)
         );
  IVDA U181 ( .A(n977), .Y(n121), .Z(n148) );
  AO2P U182 ( .A(\rem_74_2/u_div/SumTmp[1][1][6] ), .B(n628), .C(n122), .D(
        n246), .Z(n591) );
  MUX21H U183 ( .A(\rem_74_2/u_div/SumTmp[3][1][6] ), .B(
        \rem_74_2/u_div/SumTmp[7][1][6] ), .S(n103), .Z(n122) );
  AO2P U184 ( .A(n685), .B(n684), .C(n683), .D(n682), .Z(n687) );
  IVAP U185 ( .A(n757), .Z(n237) );
  B4IP U186 ( .A(n432), .Z(n429) );
  IVAP U187 ( .A(\rem_74_2/u_div/CryOut[2][0] ), .Z(n899) );
  AO7P U188 ( .A(n558), .B(n303), .C(n556), .Z(n559) );
  B2I U189 ( .A(n557), .Z2(n303) );
  IVA U190 ( .A(\rem_74_2/quotient[5] ), .Z(n308) );
  AO7P U191 ( .A(n554), .B(n303), .C(n553), .Z(n555) );
  B5I U192 ( .A(n167), .Z(n168) );
  AN2P U193 ( .A(n399), .B(n307), .Z(n301) );
  IVDA U194 ( .A(\rem_74/u_div/BInv[6][11] ), .Z(n125) );
  IV U195 ( .A(n313), .Z(n126) );
  IVAP U196 ( .A(n916), .Z(n812) );
  IVDA U197 ( .A(\rem_74/u_div/BInv[5][10] ), .Z(n127) );
  ND2P U198 ( .A(n671), .B(n670), .Z(n171) );
  IVP U199 ( .A(n356), .Z(n311) );
  B3I U200 ( .A(n292), .Z1(n357), .Z2(n358) );
  B4I U201 ( .A(n426), .Z(n424) );
  MUX21H U202 ( .A(\rem_74_2/u_div/SumTmp[2][1][6] ), .B(
        \rem_74_2/u_div/SumTmp[6][1][6] ), .S(n103), .Z(n128) );
  ND3 U203 ( .A(n551), .B(n550), .C(n549), .Z(n129) );
  ND3 U204 ( .A(n551), .B(n550), .C(n549), .Z(n552) );
  IVA U205 ( .A(n757), .Z(n130) );
  IVA U206 ( .A(n389), .Z(n391) );
  IVAP U207 ( .A(n917), .Z(n813) );
  IV U208 ( .A(n907), .Z(n853) );
  AO2P U209 ( .A(n304), .B(input_no[6]), .C(\rem_74_2/u_div/SumTmp[4][2][0] ), 
        .D(n301), .Z(n556) );
  AO2P U210 ( .A(\rem_74_2/u_div/SumTmp[1][2][0] ), .B(n304), .C(
        \rem_74_2/u_div/SumTmp[5][2][0] ), .D(n301), .Z(n553) );
  ND2 U211 ( .A(n110), .B(\rem_74_2/quotient[2] ), .Z(n898) );
  AO1P U212 ( .A(n152), .B(\rem_74/u_div/SumTmp[4][0][9] ), .C(n799), .D(n798), 
        .Z(n800) );
  ND2 U213 ( .A(n777), .B(n163), .Z(n131) );
  B5I U214 ( .A(n131), .Z(n342) );
  IVP U215 ( .A(\rem_74/u_div/CryOut[2][0] ), .Z(n777) );
  ND4P U216 ( .A(n813), .B(n812), .C(n811), .D(n336), .Z(n836) );
  OR2P U217 ( .A(\rem_74/u_div/CryOut[5][2] ), .B(n328), .Z(n671) );
  ND4P U218 ( .A(n858), .B(n857), .C(n859), .D(n856), .Z(n865) );
  IVA U219 ( .A(\rem_74_2/u_div/SumTmp[1][0][7] ), .Z(n857) );
  ND2 U220 ( .A(n881), .B(n880), .Z(n882) );
  OR2P U221 ( .A(\rem_74/u_div/CryOut[5][2] ), .B(n328), .Z(n177) );
  ND3 U222 ( .A(n132), .B(n109), .C(\rem_74_2/quotient[2] ), .Z(n902) );
  IV U223 ( .A(\rem_74_2/u_div/SumTmp[6][0][8] ), .Z(n132) );
  ND6 U224 ( .A(n133), .B(n134), .C(n135), .D(n136), .E(n137), .F(n109), .Z(
        n895) );
  IVA U225 ( .A(\rem_74_2/u_div/SumTmp[6][0][9] ), .Z(n133) );
  IVP U226 ( .A(\rem_74_2/u_div/SumTmp[6][0][2] ), .Z(n134) );
  IVP U227 ( .A(\rem_74_2/u_div/SumTmp[6][0][3] ), .Z(n135) );
  IVP U228 ( .A(\rem_74_2/u_div/SumTmp[6][0][4] ), .Z(n136) );
  IVP U229 ( .A(\rem_74_2/u_div/SumTmp[6][0][5] ), .Z(n137) );
  ND2 U230 ( .A(n651), .B(n652), .Z(n138) );
  IVAP U231 ( .A(n138), .Z(n349) );
  ND2 U232 ( .A(n648), .B(n649), .Z(n139) );
  IVAP U233 ( .A(n139), .Z(n348) );
  ND3P U234 ( .A(n140), .B(n97), .C(n141), .Z(n287) );
  IV U235 ( .A(n704), .Z(n140) );
  IVDAP U236 ( .A(n750), .Y(n937), .Z(n323) );
  AO6P U237 ( .A(\rem_74/u_div/SumTmp[4][1][8] ), .B(n173), .C(n698), .Z(n705)
         );
  EOP U238 ( .A(n509), .B(n77), .Z(n142) );
  OR2P U239 ( .A(n502), .B(n93), .Z(n509) );
  IV U240 ( .A(n505), .Z(n143) );
  IV U241 ( .A(n505), .Z(n144) );
  B5I U242 ( .A(n145), .Z(n146) );
  AN2P U243 ( .A(n613), .B(n612), .Z(n147) );
  MUX21LP U244 ( .A(n806), .B(n805), .S(n830), .Z(n916) );
  MUX21LP U245 ( .A(n796), .B(n795), .S(n830), .Z(n917) );
  IVP U246 ( .A(n736), .Z(n316) );
  OR2P U247 ( .A(n163), .B(\rem_74/u_div/CryOut[6][0] ), .Z(n149) );
  IV U248 ( .A(n773), .Z(n151) );
  IV U249 ( .A(n149), .Z(n153) );
  IV U250 ( .A(n150), .Z(n155) );
  IV U251 ( .A(n150), .Z(n156) );
  IVAP U252 ( .A(n293), .Z(n422) );
  IV U253 ( .A(n750), .Z(n157) );
  NR2 U254 ( .A(n725), .B(n769), .Z(n726) );
  B4IP U255 ( .A(n92), .Z(n255) );
  EOP U256 ( .A(n509), .B(n77), .Z(n159) );
  EOP U257 ( .A(n509), .B(n77), .Z(n160) );
  IV U258 ( .A(n293), .Z(n423) );
  IV U259 ( .A(n426), .Z(n161) );
  IVDAP U260 ( .A(n244), .Y(n145), .Z(n402) );
  IVDAP U261 ( .A(\rem_74/quotient[2] ), .Y(n163), .Z(n162) );
  B2I U262 ( .A(n292), .Z1(n158), .Z2(n164) );
  IV U263 ( .A(n759), .Z(n165) );
  IV U264 ( .A(n759), .Z(n936) );
  MUX21L U265 ( .A(\rem_74/u_div/SumTmp[6][0][0] ), .B(
        \rem_74/u_div/SumTmp[2][0][0] ), .S(n312), .Z(n803) );
  EOP U266 ( .A(n503), .B(n383), .Z(n166) );
  IVA U267 ( .A(n918), .Z(n834) );
  IVA U268 ( .A(n921), .Z(n811) );
  B5I U269 ( .A(n312), .Z(n298) );
  IVDAP U270 ( .A(n753), .Y(n172), .Z(n180) );
  ND2 U271 ( .A(n334), .B(n363), .Z(n169) );
  AN2 U272 ( .A(\rem_74/u_div/CryOut[6][2] ), .B(n240), .Z(n335) );
  IVDAP U273 ( .A(\rem_74/u_div/CryOut[6][2] ), .Y(n225), .Z(n224) );
  AN2P U274 ( .A(n66), .B(n283), .Z(n173) );
  ND3P U275 ( .A(n177), .B(n179), .C(n672), .Z(n655) );
  IVP U276 ( .A(n398), .Z(n176) );
  B4I U277 ( .A(n193), .Z(n178) );
  OR2P U278 ( .A(\rem_74/u_div/CryOut[1][2] ), .B(n221), .Z(n179) );
  IV U279 ( .A(i[2]), .Z(n181) );
  IVAP U280 ( .A(i[2]), .Z(n389) );
  ND3 U281 ( .A(i[3]), .B(i[2]), .C(i[1]), .Z(n502) );
  MUX21LP U282 ( .A(n182), .B(n183), .S(n95), .Z(n946) );
  AN2 U283 ( .A(n643), .B(n642), .Z(n182) );
  AN2 U284 ( .A(n646), .B(n645), .Z(n183) );
  MUX21LP U285 ( .A(n184), .B(n185), .S(n567), .Z(n972) );
  AN2 U286 ( .A(n513), .B(n512), .Z(n184) );
  AN2 U287 ( .A(n516), .B(n515), .Z(n185) );
  B2I U288 ( .A(n113), .Z2(n419) );
  B2I U289 ( .A(n113), .Z1(n288), .Z2(n418) );
  IVDAP U290 ( .A(n79), .Y(n83), .Z(n212) );
  B2I U291 ( .A(\rem_74_2/u_div/BInv[5][12] ), .Z2(n188) );
  AN2P U292 ( .A(n518), .B(n78), .Z(n189) );
  AN2 U293 ( .A(n399), .B(n307), .Z(n190) );
  ND3 U294 ( .A(n191), .B(n119), .C(\rem_74_2/u_div/CryOut[2][0] ), .Z(n900)
         );
  B5I U295 ( .A(i[1]), .Z(n192) );
  IVAP U296 ( .A(i[1]), .Z(n428) );
  B3IP U297 ( .A(\rem_74/quotient[8] ), .Z1(n241), .Z2(n240) );
  IV U298 ( .A(n504), .Z(n194) );
  IV U299 ( .A(n381), .Z(n382) );
  EOP U300 ( .A(n84), .B(n390), .Z(n976) );
  AN2 U301 ( .A(\rem_74/u_div/CryOut[3][2] ), .B(\rem_74/u_div/CryOut[2][2] ), 
        .Z(n205) );
  OR2P U302 ( .A(n388), .B(n506), .Z(n198) );
  IV U303 ( .A(n84), .Z(n199) );
  B2I U304 ( .A(n951), .Z2(n372) );
  MUX21LP U305 ( .A(n98), .B(n252), .S(n321), .Z(n202) );
  MUX21LP U306 ( .A(n98), .B(n252), .S(n321), .Z(n203) );
  IV U307 ( .A(i[9]), .Z(n204) );
  AO2P U308 ( .A(n335), .B(\rem_74/u_div/CryOut[7][2] ), .C(n280), .D(n205), 
        .Z(n334) );
  MUX21LP U309 ( .A(n583), .B(n582), .S(n107), .Z(n206) );
  AO11P U310 ( .A(\rem_74_2/u_div/SumTmp[1][1][8] ), .B(n105), .C(n570), .D(
        n246), .E(\rem_74_2/u_div/SumTmp[5][1][8] ), .F(n338), .Z(n583) );
  NR2 U311 ( .A(n871), .B(n870), .Z(n887) );
  IV U312 ( .A(n660), .Z(n216) );
  B5I U313 ( .A(n207), .Z(n208) );
  IV U314 ( .A(n667), .Z(n942) );
  IV U315 ( .A(n771), .Z(n209) );
  AN2P U316 ( .A(n692), .B(n691), .Z(n210) );
  AN2P U317 ( .A(n692), .B(n691), .Z(n211) );
  IVA U318 ( .A(\rem_74/u_div/SumTmp[3][0][8] ), .Z(n272) );
  AN2P U319 ( .A(n692), .B(n299), .Z(n213) );
  AN2P U320 ( .A(n692), .B(n691), .Z(n214) );
  MUX21L U321 ( .A(n272), .B(n273), .S(n315), .Z(n818) );
  MUX21L U322 ( .A(n817), .B(n816), .S(n286), .Z(n918) );
  IVAP U323 ( .A(\rem_74_2/u_div/CryOut[6][1] ), .Z(n217) );
  IV U324 ( .A(\rem_74_2/u_div/CryOut[6][1] ), .Z(n577) );
  IV U325 ( .A(\rem_74_2/u_div/CryOut[2][1] ), .Z(n249) );
  B3IP U326 ( .A(i[3]), .Z1(n384), .Z2(n383) );
  NR2P U327 ( .A(n219), .B(n632), .Z(n633) );
  IVDA U328 ( .A(n329), .Z(n300) );
  OR2 U329 ( .A(n508), .B(n264), .Z(n220) );
  OR3P U330 ( .A(n499), .B(n387), .C(n497), .Z(n508) );
  IV U331 ( .A(\rem_74_2/u_div/BInv[6][13] ), .Z(n222) );
  IVA U332 ( .A(n222), .Z(n223) );
  ENP U333 ( .A(n509), .B(n77), .Z(n350) );
  IV U334 ( .A(n309), .Z(n310) );
  IVAP U335 ( .A(n258), .Z(n268) );
  EOP U336 ( .A(n368), .B(n360), .Z(n226) );
  IV U337 ( .A(n629), .Z(n227) );
  IVA U338 ( .A(n628), .Z(n228) );
  AO2P U339 ( .A(n763), .B(n762), .C(n761), .D(n760), .Z(n770) );
  IVDA U340 ( .A(n769), .Y(n230), .Z(n229) );
  IVDAP U341 ( .A(\rem_74_2/u_div/CryOut[6][2] ), .Y(n307), .Z(n306) );
  MUX21LP U342 ( .A(n345), .B(n344), .S(n637), .Z(n956) );
  IVP U343 ( .A(n231), .Z(n232) );
  IVP U344 ( .A(\rem_74/u_div/SumTmp[7][0][8] ), .Z(n273) );
  IVDAP U345 ( .A(n978), .Y(n231), .Z(n414) );
  ND4 U346 ( .A(n353), .B(n500), .C(n285), .D(n427), .Z(n501) );
  IVDAP U347 ( .A(n241), .Y(n233), .Z(n280) );
  MUX21L U348 ( .A(n821), .B(n820), .S(n830), .Z(n920) );
  MUX21LP U349 ( .A(n589), .B(n588), .S(n107), .Z(
        \rem_74_2/u_div/PartRem[1][10] ) );
  B2I U350 ( .A(\rem_74/u_div/CryOut[7][1] ), .Z2(n234) );
  B5I U351 ( .A(i[8]), .Z(n261) );
  MUX21LP U352 ( .A(n620), .B(n619), .S(n147), .Z(n236) );
  AO11P U353 ( .A(\rem_74_2/u_div/SumTmp[5][1][2] ), .B(n338), .C(
        \rem_74_2/u_div/SumTmp[1][1][2] ), .D(n628), .E(n246), .F(n616), .Z(
        n620) );
  ND2P U354 ( .A(i[5]), .B(i[4]), .Z(n497) );
  IVA U355 ( .A(n940), .Z(n238) );
  IVP U356 ( .A(n238), .Z(n239) );
  IVDA U357 ( .A(\rem_74/u_div/BInv[7][9] ), .Z(n242) );
  B2IP U358 ( .A(n374), .Z1(n398), .Z2(n386) );
  B2I U359 ( .A(\rem_74/u_div/BInv[6][6] ), .Z2(n243) );
  EOP U360 ( .A(n508), .B(n92), .Z(n244) );
  B5I U361 ( .A(n505), .Z(n974) );
  AO6P U362 ( .A(\rem_74_2/u_div/SumTmp[4][1][1] ), .B(n338), .C(n624), .Z(
        n625) );
  B4IP U363 ( .A(n428), .Z(n427) );
  IVAP U364 ( .A(n601), .Z(n635) );
  IVAP U365 ( .A(n597), .Z(n636) );
  IVDA U366 ( .A(\rem_74/u_div/BInv[6][10] ), .Z(n245) );
  MUX21L U367 ( .A(n810), .B(n809), .S(n286), .Z(n921) );
  MUX21LP U368 ( .A(n108), .B(n71), .S(n107), .Z(n960) );
  AN2P U369 ( .A(n591), .B(n590), .Z(n247) );
  IVA U370 ( .A(n169), .Z(n248) );
  B3IP U371 ( .A(n630), .Z1(n246), .Z2(n295) );
  B5IP U372 ( .A(n319), .Z(n338) );
  IVAP U373 ( .A(\rem_74_2/u_div/CryOut[2][1] ), .Z(n578) );
  EOP U374 ( .A(n507), .B(n385), .Z(n250) );
  B4IP U375 ( .A(n250), .Z(n362) );
  B4IP U376 ( .A(n268), .Z(n271) );
  B2IP U377 ( .A(n978), .Z1(n75), .Z2(n413) );
  AO4P U378 ( .A(n287), .B(n749), .C(n74), .D(n748), .Z(n750) );
  IVA U379 ( .A(n782), .Z(n830) );
  IVAP U380 ( .A(n782), .Z(n286) );
  IVDA U381 ( .A(n242), .Z(n251) );
  IVAP U382 ( .A(i[8]), .Z(n950) );
  NR3P U383 ( .A(n199), .B(n284), .C(n498), .Z(n368) );
  IV U384 ( .A(n827), .Z(n253) );
  IVAP U385 ( .A(n92), .Z(n254) );
  IVDA U386 ( .A(\rem_74/u_div/BInv[3][2] ), .Z(n256) );
  IV U387 ( .A(n759), .Z(n257) );
  EOP U388 ( .A(n502), .B(n94), .Z(n258) );
  B2IP U389 ( .A(n244), .Z2(n401) );
  AO6P U390 ( .A(\rem_74_2/u_div/SumTmp[4][1][2] ), .B(n338), .C(n618), .Z(
        n619) );
  ND2P U391 ( .A(\rem_74_2/u_div/CryOut[5][1] ), .B(n217), .Z(n575) );
  IVDA U392 ( .A(\rem_74/u_div/BInv[7][5] ), .Z(n259) );
  EOP U393 ( .A(n508), .B(n92), .Z(n980) );
  IVDA U394 ( .A(\rem_74_2/u_div/BInv[3][10] ), .Z(n260) );
  IVA U395 ( .A(\rem_74_2/u_div/CryOut[3][1] ), .Z(n278) );
  ND2P U396 ( .A(\rem_74/u_div/SumTmp[1][3][1] ), .B(
        \rem_74/u_div/CryOut[1][3] ), .Z(n639) );
  B2IP U397 ( .A(n951), .Z1(n201), .Z2(n371) );
  IVDA U398 ( .A(n245), .Z(n262) );
  IVA U399 ( .A(n941), .Z(n322) );
  B2I U400 ( .A(\rem_74/u_div/BInv[3][5] ), .Z2(n263) );
  ND3 U401 ( .A(n353), .B(i[8]), .C(n120), .Z(n264) );
  AN2 U402 ( .A(i[7]), .B(i[6]), .Z(n353) );
  ND4P U403 ( .A(n354), .B(n285), .C(n382), .D(n427), .Z(n507) );
  ND3 U404 ( .A(\rem_74/u_div/CryOut[5][0] ), .B(n162), .C(n69), .Z(n778) );
  B5I U405 ( .A(n266), .Z(n267) );
  OR2P U406 ( .A(n163), .B(\rem_74/u_div/CryOut[6][0] ), .Z(n773) );
  IVAP U407 ( .A(n268), .Z(n270) );
  MUX21LP U408 ( .A(input_no[9]), .B(\rem_74_2/u_div/SumTmp[1][3][0] ), .S(
        \rem_74_2/u_div/CryOut[1][3] ), .Z(n510) );
  B4IP U409 ( .A(n510), .Z(n973) );
  MUX21L U410 ( .A(n274), .B(n275), .S(n315), .Z(n814) );
  MUX21L U411 ( .A(n276), .B(n277), .S(n315), .Z(n807) );
  B2IP U412 ( .A(n374), .Z1(n193), .Z2(n411) );
  MUX21LP U413 ( .A(n348), .B(n349), .S(n248), .Z(n333) );
  MUX21LP U414 ( .A(n348), .B(n349), .S(n248), .Z(n332) );
  MUX21LP U415 ( .A(n348), .B(n349), .S(n248), .Z(n945) );
  B2I U416 ( .A(n979), .Z2(n400) );
  B4I U417 ( .A(n78), .Z(n399) );
  B2IP U418 ( .A(n933), .Z1(n266), .Z2(n281) );
  B3I U419 ( .A(n114), .Z1(n285), .Z2(n284) );
  AO4P U420 ( .A(n770), .B(n229), .C(n230), .D(n768), .Z(n771) );
  ND3 U421 ( .A(n79), .B(n307), .C(\rem_74_2/u_div/CryOut[5][2] ), .Z(n549) );
  IV U422 ( .A(n766), .Z(n764) );
  MUX21LP U423 ( .A(n713), .B(n712), .S(n237), .Z(
        \rem_74/u_div/PartRem[1][10] ) );
  MUX21LP U424 ( .A(n706), .B(n705), .S(n237), .Z(
        \rem_74/u_div/PartRem[1][11] ) );
  AO4P U425 ( .A(n287), .B(n735), .C(n74), .D(n734), .Z(n736) );
  IVP U426 ( .A(n576), .Z(n613) );
  MUX21LP U427 ( .A(n294), .B(n282), .S(n293), .Z(n769) );
  AO3P U428 ( .A(n781), .B(n780), .C(n779), .D(n778), .Z(n782) );
  MUX21LP U429 ( .A(n636), .B(n635), .S(n107), .Z(n959) );
  ND2P U430 ( .A(n792), .B(n791), .Z(n923) );
  AO4 U431 ( .A(n928), .B(n929), .C(n289), .D(\state[0] ), .Z(n934) );
  B2I U432 ( .A(n270), .Z2(n290) );
  MUX21LP U433 ( .A(n566), .B(n565), .S(n562), .Z(n964) );
  IVAP U434 ( .A(n548), .Z(n565) );
  AO2P U435 ( .A(n292), .B(n701), .C(n700), .D(n65), .Z(n702) );
  ND2P U436 ( .A(\rem_74/u_div/CryOut[3][1] ), .B(\rem_74/u_div/CryOut[2][1] ), 
        .Z(n700) );
  B3I U437 ( .A(n667), .Z1(n291), .Z2(n207) );
  B3IP U438 ( .A(\rem_74/quotient[5] ), .Z1(n293), .Z2(n292) );
  ND2P U439 ( .A(\rem_74/u_div/CryOut[5][1] ), .B(n699), .Z(n701) );
  ND2P U440 ( .A(\rem_74_2/u_div/CryOut[1][1] ), .B(n578), .Z(n574) );
  AN2 U441 ( .A(n177), .B(n179), .Z(n296) );
  NR2P U442 ( .A(n887), .B(n886), .Z(n888) );
  ND2P U443 ( .A(n885), .B(n884), .Z(n886) );
  MUX21LP U444 ( .A(\rem_74/u_div/CryOut[3][2] ), .B(
        \rem_74/u_div/CryOut[7][2] ), .S(n233), .Z(n682) );
  B3IP U445 ( .A(\rem_74/quotient[2] ), .Z1(n312), .Z2(n315) );
  MUX21LP U446 ( .A(n583), .B(n582), .S(n107), .Z(
        \rem_74_2/u_div/PartRem[1][11] ) );
  OR2 U447 ( .A(n679), .B(n678), .Z(n691) );
  MUX21LP U448 ( .A(n247), .B(n71), .S(n107), .Z(n961) );
  EOP U449 ( .A(n220), .B(n100), .Z(n977) );
  MUX21LP U450 ( .A(n564), .B(n563), .S(n567), .Z(n966) );
  MUX21LP U451 ( .A(n561), .B(n560), .S(n567), .Z(n970) );
  IVAP U452 ( .A(n129), .Z(n562) );
  OR2P U453 ( .A(n673), .B(n674), .Z(n692) );
  AN2P U454 ( .A(n79), .B(n307), .Z(n302) );
  B2I U455 ( .A(n80), .Z1(n365), .Z2(n404) );
  AN2P U456 ( .A(n518), .B(n83), .Z(n305) );
  MUX21LP U457 ( .A(n306), .B(\rem_74_2/u_div/CryOut[2][2] ), .S(n78), .Z(n557) );
  IV U458 ( .A(\rem_74_2/u_div/CryOut[2][2] ), .Z(n518) );
  MUX21H U459 ( .A(\rem_74/u_div/CryOut[2][2] ), .B(
        \rem_74/u_div/CryOut[6][2] ), .S(n240), .Z(n309) );
  AO4P U460 ( .A(n424), .B(n578), .C(n308), .D(n577), .Z(n580) );
  MUX21LP U461 ( .A(n569), .B(n568), .S(n567), .Z(n962) );
  IVAP U462 ( .A(n552), .Z(n567) );
  IV U463 ( .A(n736), .Z(n317) );
  IV U464 ( .A(n736), .Z(n939) );
  MUX21LP U465 ( .A(n743), .B(n742), .S(n130), .Z(n318) );
  B4IP U466 ( .A(n318), .Z(n938) );
  OR2P U467 ( .A(n308), .B(\rem_74_2/u_div/CryOut[6][1] ), .Z(n319) );
  IV U468 ( .A(n119), .Z(n320) );
  IV U469 ( .A(\rem_74/u_div/CryOut[1][3] ), .Z(n321) );
  ND4P U470 ( .A(n834), .B(n833), .C(n341), .D(n346), .Z(n835) );
  ND2P U471 ( .A(n613), .B(n612), .Z(n581) );
  ND2P U472 ( .A(n580), .B(n579), .Z(n612) );
  B5I U473 ( .A(n323), .Z(n324) );
  AO3P U474 ( .A(n891), .B(n890), .C(n889), .D(n888), .Z(n915) );
  MUX21LP U475 ( .A(\rem_74_2/u_div/CryOut[6][1] ), .B(
        \rem_74_2/u_div/CryOut[2][1] ), .S(n426), .Z(n630) );
  NR2P U476 ( .A(n929), .B(n928), .Z(n930) );
  ND2P U477 ( .A(n892), .B(n915), .Z(n928) );
  ND2 U478 ( .A(n463), .B(n327), .Z(n325) );
  AN2 U479 ( .A(n325), .B(n326), .Z(n465) );
  OR2 U480 ( .A(n932), .B(n464), .Z(n326) );
  AN2P U481 ( .A(n462), .B(\state[0] ), .Z(n327) );
  OR2P U482 ( .A(n388), .B(n506), .Z(n329) );
  OR2P U483 ( .A(n388), .B(n506), .Z(n330) );
  IVP U484 ( .A(n167), .Z(n331) );
  B2I U485 ( .A(n166), .Z2(n417) );
  AO6 U486 ( .A(n869), .B(n868), .C(n119), .Z(n870) );
  ND2 U487 ( .A(\rem_74_2/u_div/CryOut[1][0] ), .B(n899), .Z(n867) );
  B2IP U488 ( .A(n166), .Z2(n415) );
  IV U489 ( .A(\rem_74_2/u_div/SumTmp[7][0][9] ), .Z(n846) );
  IV U490 ( .A(\rem_74_2/u_div/SumTmp[7][0][7] ), .Z(n848) );
  IV U491 ( .A(\rem_74_2/u_div/SumTmp[7][0][8] ), .Z(n847) );
  IVAP U492 ( .A(n686), .Z(n676) );
  AO7P U493 ( .A(n877), .B(n876), .C(n86), .Z(n885) );
  ND2P U494 ( .A(n875), .B(n874), .Z(n876) );
  IV U495 ( .A(\rem_74_2/u_div/SumTmp[5][0][4] ), .Z(n873) );
  AO7P U496 ( .A(n883), .B(n882), .C(n96), .Z(n884) );
  IV U497 ( .A(\rem_74_2/u_div/SumTmp[1][0][4] ), .Z(n879) );
  MUX21H U498 ( .A(n801), .B(n800), .S(n286), .Z(n336) );
  ND2P U499 ( .A(n102), .B(n914), .Z(n929) );
  IV U500 ( .A(n427), .Z(n430) );
  AO4P U501 ( .A(n903), .B(n902), .C(n901), .D(n900), .Z(n904) );
  IVP U502 ( .A(n94), .Z(n351) );
  B2I U503 ( .A(n87), .Z2(n409) );
  AN2 U504 ( .A(n442), .B(n441), .Z(n337) );
  MUX21LP U505 ( .A(n395), .B(n396), .S(\rem_74_2/u_div/CryOut[1][3] ), .Z(
        n394) );
  EOP U506 ( .A(n62), .B(n360), .Z(n355) );
  AN2 U507 ( .A(i[5]), .B(i[4]), .Z(n354) );
  ND2 U508 ( .A(\rem_74_2/u_div/CryOut[5][0] ), .B(n110), .Z(n869) );
  AN2P U509 ( .A(n422), .B(n283), .Z(n339) );
  AN2P U510 ( .A(n613), .B(n612), .Z(n340) );
  MUX21L U511 ( .A(n784), .B(n783), .S(n286), .Z(n792) );
  MUX21L U512 ( .A(n790), .B(n789), .S(n286), .Z(n791) );
  IVP U513 ( .A(\rem_74_2/u_div/SumTmp[5][0][9] ), .Z(n874) );
  IVP U514 ( .A(\rem_74_2/u_div/SumTmp[5][0][8] ), .Z(n875) );
  MUX21H U515 ( .A(n825), .B(n824), .S(n286), .Z(n341) );
  AO6 U516 ( .A(\rem_74_2/u_div/SumTmp[4][1][8] ), .B(n338), .C(n573), .Z(n582) );
  IVP U517 ( .A(\rem_74_2/u_div/SumTmp[3][0][9] ), .Z(n837) );
  ND4 U518 ( .A(n839), .B(n838), .C(n73), .D(n837), .Z(n845) );
  IVP U519 ( .A(\rem_74_2/u_div/SumTmp[3][0][7] ), .Z(n839) );
  IVP U520 ( .A(\rem_74_2/u_div/SumTmp[3][0][8] ), .Z(n838) );
  IVP U521 ( .A(\rem_74_2/u_div/SumTmp[1][0][6] ), .Z(n878) );
  IVP U522 ( .A(\rem_74_2/u_div/SumTmp[5][0][6] ), .Z(n872) );
  NR2 U523 ( .A(n680), .B(n171), .Z(n689) );
  ND2 U524 ( .A(\rem_74_2/u_div/CryOut[3][0] ), .B(
        \rem_74_2/u_div/CryOut[2][0] ), .Z(n866) );
  AN2P U525 ( .A(n265), .B(n225), .Z(n343) );
  IVP U526 ( .A(\rem_74_2/u_div/SumTmp[5][0][7] ), .Z(n861) );
  AN2P U527 ( .A(n607), .B(n606), .Z(n344) );
  AN2P U528 ( .A(n604), .B(n603), .Z(n345) );
  IVP U529 ( .A(\rem_74_2/u_div/SumTmp[1][0][9] ), .Z(n880) );
  IVP U530 ( .A(\rem_74_2/u_div/SumTmp[1][0][8] ), .Z(n881) );
  MUX21H U531 ( .A(n832), .B(n831), .S(n286), .Z(n346) );
  AO6 U532 ( .A(\rem_74_2/u_div/SumTmp[4][1][7] ), .B(n338), .C(n587), .Z(n588) );
  NR2 U533 ( .A(n845), .B(n844), .Z(n891) );
  AO2 U534 ( .A(n96), .B(n865), .C(n86), .D(n864), .Z(n889) );
  AO7 U535 ( .A(n296), .B(n681), .C(n686), .Z(n688) );
  AN2P U536 ( .A(n529), .B(n528), .Z(n347) );
  NR2 U537 ( .A(\rem_74_2/u_div/SumTmp[3][0][5] ), .B(
        \rem_74_2/u_div/SumTmp[3][0][6] ), .Z(n842) );
  NR2 U538 ( .A(\rem_74_2/u_div/SumTmp[7][0][5] ), .B(
        \rem_74_2/u_div/SumTmp[7][0][6] ), .Z(n851) );
  MUX21L U539 ( .A(n480), .B(n479), .S(n378), .Z(n986) );
  ND4 U540 ( .A(n863), .B(n862), .C(n861), .D(n860), .Z(n864) );
  IVP U541 ( .A(\rem_74_2/u_div/SumTmp[5][0][0] ), .Z(n862) );
  NR2 U542 ( .A(\rem_74_2/u_div/SumTmp[5][0][3] ), .B(
        \rem_74_2/u_div/SumTmp[5][0][2] ), .Z(n863) );
  NR2 U543 ( .A(\rem_74_2/u_div/SumTmp[5][0][5] ), .B(
        \rem_74_2/u_div/SumTmp[5][0][1] ), .Z(n860) );
  IVP U544 ( .A(\rem_74_2/u_div/SumTmp[1][0][0] ), .Z(n858) );
  NR2 U545 ( .A(\rem_74_2/u_div/SumTmp[1][0][3] ), .B(
        \rem_74_2/u_div/SumTmp[1][0][2] ), .Z(n859) );
  NR2 U546 ( .A(\rem_74_2/u_div/SumTmp[1][0][5] ), .B(
        \rem_74_2/u_div/SumTmp[1][0][1] ), .Z(n856) );
  AN2P U547 ( .A(n532), .B(n531), .Z(n352) );
  AO6 U548 ( .A(\rem_74/u_div/SumTmp[4][1][7] ), .B(n173), .C(n711), .Z(n712)
         );
  ND4 U549 ( .A(n843), .B(n842), .C(n841), .D(n840), .Z(n844) );
  IVP U550 ( .A(\rem_74_2/u_div/SumTmp[3][0][2] ), .Z(n841) );
  NR2 U551 ( .A(\rem_74_2/u_div/SumTmp[3][0][1] ), .B(
        \rem_74_2/u_div/SumTmp[3][0][3] ), .Z(n843) );
  NR2 U552 ( .A(\rem_74_2/u_div/SumTmp[3][0][0] ), .B(
        \rem_74_2/u_div/SumTmp[3][0][4] ), .Z(n840) );
  ND4 U553 ( .A(n852), .B(n851), .C(n850), .D(n849), .Z(n854) );
  IVP U554 ( .A(\rem_74_2/u_div/SumTmp[7][0][2] ), .Z(n850) );
  NR2 U555 ( .A(\rem_74_2/u_div/SumTmp[7][0][1] ), .B(
        \rem_74_2/u_div/SumTmp[7][0][3] ), .Z(n852) );
  NR2 U556 ( .A(\rem_74_2/u_div/SumTmp[7][0][0] ), .B(
        \rem_74_2/u_div/SumTmp[7][0][4] ), .Z(n849) );
  AO7 U557 ( .A(N41), .B(n434), .C(n452), .Z(n444) );
  AO6 U558 ( .A(n494), .B(n466), .C(n484), .Z(n481) );
  AO6 U559 ( .A(N44), .B(n640), .C(N45), .Z(n461) );
  EO U560 ( .A(n419), .B(n474), .Z(n477) );
  IVA U561 ( .A(input_no[9]), .Z(n395) );
  IVA U562 ( .A(\rem_74_2/u_div/SumTmp[1][3][0] ), .Z(n396) );
  MUX21L U563 ( .A(n490), .B(n491), .S(n89), .Z(n991) );
  IVP U564 ( .A(input_no[5]), .Z(n982) );
  AO6 U565 ( .A(is_prime), .B(n102), .C(n919), .Z(n925) );
  IV U566 ( .A(n963), .Z(n609) );
  AN2 U567 ( .A(\rem_74/u_div/SumTmp[2][0][9] ), .B(n67), .Z(n798) );
  B2IP U568 ( .A(n292), .Z1(n356), .Z2(n359) );
  B4IP U569 ( .A(\rem_74_2/quotient[5] ), .Z(n426) );
  B4IP U570 ( .A(i[9]), .Z(n360) );
  ND2 U571 ( .A(\rem_74/u_div/SumTmp[1][3][2] ), .B(
        \rem_74/u_div/CryOut[1][3] ), .Z(n638) );
  ND3 U572 ( .A(n177), .B(n179), .C(n672), .Z(n363) );
  OR2P U573 ( .A(\rem_74/u_div/CryOut[1][2] ), .B(n221), .Z(n670) );
  AN2P U574 ( .A(n686), .B(n280), .Z(n364) );
  EOP U575 ( .A(n507), .B(n201), .Z(n979) );
  AO4P U576 ( .A(n682), .B(n672), .C(n309), .D(n171), .Z(n674) );
  ND2P U577 ( .A(reset_n), .B(n465), .Z(n484) );
  ND2P U578 ( .A(n475), .B(\state[0] ), .Z(n476) );
  B5I U579 ( .A(n484), .Z(n475) );
  EOP U580 ( .A(n501), .B(n380), .Z(n978) );
  IVAP U581 ( .A(n497), .Z(n500) );
  IVAP U582 ( .A(i[7]), .Z(n951) );
  AO6 U583 ( .A(n494), .B(n469), .C(n484), .Z(n479) );
  AO6 U584 ( .A(n494), .B(n360), .C(n493), .Z(n495) );
  B2I U585 ( .A(n374), .Z1(n373), .Z2(n410) );
  MUX21LP U586 ( .A(n561), .B(n560), .S(n567), .Z(n971) );
  MUX21LP U587 ( .A(n564), .B(n563), .S(n562), .Z(n967) );
  AO2P U588 ( .A(n424), .B(n575), .C(n574), .D(n308), .Z(n576) );
  MUX21LP U589 ( .A(n347), .B(n352), .S(n562), .Z(n968) );
  ND2P U590 ( .A(\rem_74_2/u_div/SumTmp[1][3][2] ), .B(
        \rem_74_2/u_div/CryOut[1][3] ), .Z(n504) );
  AO3 U591 ( .A(\rem_74_2/u_div/CryOut[3][2] ), .B(n518), .C(n517), .D(n78), 
        .Z(n551) );
  ND4 U592 ( .A(n848), .B(n847), .C(n320), .D(n846), .Z(n855) );
  AO6 U593 ( .A(n867), .B(n866), .C(n72), .Z(n871) );
  EOP U594 ( .A(n220), .B(n100), .Z(n933) );
  NR2 U595 ( .A(n722), .B(n753), .Z(n724) );
  ND2P U596 ( .A(n694), .B(n693), .Z(n660) );
  AO4P U597 ( .A(n666), .B(n169), .C(n95), .D(n665), .Z(n667) );
  AO4P U598 ( .A(n689), .B(n688), .C(n687), .D(n686), .Z(n690) );
  IV U599 ( .A(n674), .Z(n679) );
  AO7 U600 ( .A(n741), .B(n229), .C(n740), .Z(n742) );
  AO7 U601 ( .A(n738), .B(n229), .C(n737), .Z(n743) );
  NR2 U602 ( .A(n717), .B(n769), .Z(n718) );
  NR2 U603 ( .A(n714), .B(n769), .Z(n716) );
  ND2 U604 ( .A(\rem_74_2/u_div/CryOut[7][0] ), .B(n109), .Z(n868) );
  MUX21LP U605 ( .A(n615), .B(n614), .S(n147), .Z(n955) );
  MUX21LP U606 ( .A(n634), .B(n633), .S(n340), .Z(n952) );
  AO4P U607 ( .A(n758), .B(n287), .C(n74), .D(n756), .Z(n759) );
  MUX21LP U608 ( .A(n620), .B(n619), .S(n147), .Z(n954) );
  MUX21LP U609 ( .A(n569), .B(n568), .S(n567), .Z(n963) );
  MUX21LP U610 ( .A(n345), .B(n344), .S(n637), .Z(n957) );
  NR8 U611 ( .A(\rem_74_2/u_div/SumTmp[4][0][8] ), .B(
        \rem_74_2/u_div/SumTmp[4][0][9] ), .C(n898), .D(
        \rem_74_2/u_div/CryOut[5][0] ), .E(\rem_74_2/u_div/SumTmp[4][0][6] ), 
        .F(\rem_74_2/u_div/SumTmp[4][0][3] ), .G(
        \rem_74_2/u_div/SumTmp[4][0][0] ), .H(\rem_74_2/u_div/SumTmp[4][0][4] ), .Z(n905) );
  MUX21LP U612 ( .A(n347), .B(n352), .S(n562), .Z(n969) );
  MUX21LP U613 ( .A(n626), .B(n625), .S(n340), .Z(n953) );
  MUX21L U614 ( .A(n932), .B(n931), .S(n930), .Z(n57) );
  OR3P U615 ( .A(n704), .B(n703), .C(n702), .Z(n757) );
  MUX21LP U616 ( .A(n721), .B(n720), .S(n130), .Z(n941) );
  MUX21LP U617 ( .A(n729), .B(n728), .S(n237), .Z(n940) );
  MUX21LP U618 ( .A(\rem_74/u_div/CryOut[2][2] ), .B(n224), .S(n240), .Z(n672)
         );
  AO12 U619 ( .A(n320), .B(n909), .C(n73), .D(n908), .E(n907), .F(n906), .G(
        n905), .H(n904), .Z(n914) );
  ND2P U620 ( .A(n249), .B(n426), .Z(n629) );
  MUX21LP U621 ( .A(n566), .B(n565), .S(n562), .Z(n965) );
  ND2P U622 ( .A(\rem_74_2/u_div/SumTmp[1][3][1] ), .B(
        \rem_74_2/u_div/CryOut[1][3] ), .Z(n505) );
  MUX21LP U623 ( .A(n636), .B(n635), .S(n107), .Z(n958) );
  B4IP U624 ( .A(n639), .Z(n948) );
  B5IP U625 ( .A(n350), .Z(n420) );
  B5I U626 ( .A(n476), .Z(n494) );
  B5I U627 ( .A(n629), .Z(n628) );
  MUX21LP U628 ( .A(\rem_74/u_div/CryOut[2][2] ), .B(n224), .S(n175), .Z(n686)
         );
  MUX21LP U629 ( .A(n282), .B(n294), .S(n292), .Z(n753) );
  MUX21LP U630 ( .A(\rem_74/u_div/CryOut[2][0] ), .B(
        \rem_74/u_div/CryOut[6][0] ), .S(\rem_74/quotient[2] ), .Z(n828) );
  IVA U631 ( .A(input_no[7]), .Z(n435) );
  ND2 U632 ( .A(n430), .B(n361), .Z(n474) );
  ND2 U633 ( .A(n474), .B(n288), .Z(n469) );
  IVA U634 ( .A(n469), .Z(n478) );
  ND2 U635 ( .A(n478), .B(n354), .Z(n466) );
  IVA U636 ( .A(n466), .Z(n483) );
  AN2P U637 ( .A(n483), .B(n385), .Z(n437) );
  MUX21L U638 ( .A(n200), .B(n437), .S(n92), .Z(n467) );
  OR2 U639 ( .A(N0), .B(N1), .Z(n438) );
  IVA U640 ( .A(input_no[9]), .Z(n640) );
  IVA U641 ( .A(input_no[4]), .Z(n622) );
  IVA U642 ( .A(input_no[2]), .Z(n443) );
  ND8 U643 ( .A(n640), .B(n436), .C(n435), .D(n434), .E(n982), .F(n622), .G(
        n433), .H(n443), .Z(n910) );
  ND4 U644 ( .A(input_no[0]), .B(\state[0] ), .C(n438), .D(n910), .Z(n913) );
  IVA U645 ( .A(n913), .Z(n464) );
  ND2 U646 ( .A(N42), .B(n435), .Z(n459) );
  ND2 U647 ( .A(N43), .B(n436), .Z(n458) );
  IVA U648 ( .A(N42), .Z(n439) );
  ND2 U649 ( .A(input_no[7]), .B(n439), .Z(n452) );
  IVA U650 ( .A(n444), .Z(n456) );
  IVA U651 ( .A(N40), .Z(n442) );
  IVA U652 ( .A(n982), .Z(n441) );
  ND2 U653 ( .A(N39), .B(n622), .Z(n440) );
  AO4 U654 ( .A(n442), .B(n441), .C(n337), .D(n440), .Z(n455) );
  IVA U655 ( .A(N38), .Z(n451) );
  AO2 U656 ( .A(n981), .B(N35), .C(N37), .D(n443), .Z(n445) );
  ND2 U657 ( .A(N38), .B(n433), .Z(n447) );
  AO1P U658 ( .A(n445), .B(n447), .C(n337), .D(n444), .Z(n446) );
  IVA U659 ( .A(n446), .Z(n450) );
  ND2 U660 ( .A(input_no[2]), .B(n447), .Z(n448) );
  AO4 U661 ( .A(N39), .B(n622), .C(N37), .D(n448), .Z(n449) );
  AO1P U662 ( .A(input_no[3]), .B(n451), .C(n450), .D(n449), .Z(n454) );
  AN3 U663 ( .A(N41), .B(n434), .C(n452), .Z(n453) );
  AO1P U664 ( .A(n456), .B(n455), .C(n454), .D(n453), .Z(n457) );
  ND4 U665 ( .A(n461), .B(n459), .C(n458), .D(n457), .Z(n463) );
  AO4 U666 ( .A(N44), .B(n640), .C(N43), .D(n436), .Z(n460) );
  ND2 U667 ( .A(n461), .B(n460), .Z(n462) );
  ND2 U668 ( .A(n463), .B(n462), .Z(n912) );
  AO4 U669 ( .A(n467), .B(n476), .C(n371), .D(n481), .Z(n989) );
  AN2P U670 ( .A(n478), .B(n404), .Z(n468) );
  MUX21L U671 ( .A(n365), .B(n468), .S(n377), .Z(n470) );
  AO4 U672 ( .A(n470), .B(n476), .C(n404), .D(n479), .Z(n987) );
  MUX21L U673 ( .A(n476), .B(n475), .S(n429), .Z(n984) );
  ND2 U674 ( .A(n494), .B(n409), .Z(n472) );
  MUX21L U675 ( .A(n81), .B(n932), .S(n475), .Z(n471) );
  ND2 U676 ( .A(n472), .B(n471), .Z(n59) );
  ND2 U677 ( .A(n475), .B(n932), .Z(n473) );
  ND2 U678 ( .A(n176), .B(n473), .Z(n60) );
  AO4 U679 ( .A(n477), .B(n476), .C(n418), .D(n475), .Z(n985) );
  ND2 U680 ( .A(n494), .B(n478), .Z(n480) );
  ND2 U681 ( .A(n494), .B(n483), .Z(n482) );
  MUX21L U682 ( .A(n482), .B(n481), .S(n92), .Z(n988) );
  ND2 U683 ( .A(n483), .B(n353), .Z(n485) );
  IVA U684 ( .A(n485), .Z(n487) );
  ND2 U685 ( .A(n494), .B(n487), .Z(n486) );
  AO6P U686 ( .A(n494), .B(n485), .C(n484), .Z(n489) );
  MUX21L U687 ( .A(n486), .B(n489), .S(n380), .Z(n990) );
  ND3 U688 ( .A(n487), .B(n380), .C(n494), .Z(n491) );
  ND2 U689 ( .A(n494), .B(n90), .Z(n488) );
  ND2 U690 ( .A(n489), .B(n488), .Z(n493) );
  IVA U691 ( .A(n493), .Z(n490) );
  IVA U692 ( .A(n491), .Z(n492) );
  ND2 U693 ( .A(n492), .B(n88), .Z(n496) );
  MUX21L U694 ( .A(n496), .B(n495), .S(n100), .Z(n983) );
  ND2 U695 ( .A(i[2]), .B(i[1]), .Z(n503) );
  MUX21L U696 ( .A(\rem_74_2/u_div/SumTmp[3][2][5] ), .B(
        \rem_74_2/u_div/SumTmp[7][2][5] ), .S(n399), .Z(n511) );
  EO1 U697 ( .A(\rem_74_2/u_div/SumTmp[5][2][5] ), .B(n302), .C(n557), .D(n511), .Z(n513) );
  ND2 U698 ( .A(\rem_74_2/u_div/SumTmp[1][2][5] ), .B(n305), .Z(n512) );
  MUX21L U699 ( .A(\rem_74_2/u_div/SumTmp[2][2][5] ), .B(
        \rem_74_2/u_div/SumTmp[6][2][5] ), .S(n399), .Z(n514) );
  EO1 U700 ( .A(\rem_74_2/u_div/SumTmp[4][2][5] ), .B(n302), .C(n557), .D(n514), .Z(n516) );
  ND2 U701 ( .A(n194), .B(n305), .Z(n515) );
  OR2 U702 ( .A(\rem_74_2/u_div/CryOut[1][2] ), .B(
        \rem_74_2/u_div/CryOut[2][2] ), .Z(n517) );
  ND3 U703 ( .A(n306), .B(n79), .C(\rem_74_2/u_div/CryOut[7][2] ), .Z(n550) );
  MUX21L U704 ( .A(\rem_74_2/u_div/SumTmp[3][2][4] ), .B(
        \rem_74_2/u_div/SumTmp[7][2][4] ), .S(n399), .Z(n519) );
  EO1 U705 ( .A(\rem_74_2/u_div/SumTmp[5][2][4] ), .B(n302), .C(n557), .D(n519), .Z(n521) );
  ND2 U706 ( .A(\rem_74_2/u_div/SumTmp[1][2][4] ), .B(n305), .Z(n520) );
  ND2 U707 ( .A(n521), .B(n520), .Z(n522) );
  IVA U708 ( .A(n522), .Z(n561) );
  MUX21L U709 ( .A(\rem_74_2/u_div/SumTmp[2][2][4] ), .B(
        \rem_74_2/u_div/SumTmp[6][2][4] ), .S(n399), .Z(n523) );
  EO1 U710 ( .A(\rem_74_2/u_div/SumTmp[4][2][4] ), .B(n302), .C(n557), .D(n523), .Z(n525) );
  ND2 U711 ( .A(n144), .B(n305), .Z(n524) );
  ND2 U712 ( .A(n525), .B(n524), .Z(n526) );
  IVA U713 ( .A(n526), .Z(n560) );
  MUX21L U714 ( .A(\rem_74_2/u_div/SumTmp[3][2][3] ), .B(
        \rem_74_2/u_div/SumTmp[7][2][3] ), .S(n399), .Z(n527) );
  EO1 U715 ( .A(\rem_74_2/u_div/SumTmp[5][2][3] ), .B(n190), .C(n557), .D(n527), .Z(n529) );
  ND2 U716 ( .A(\rem_74_2/u_div/SumTmp[1][2][3] ), .B(n305), .Z(n528) );
  MUX21L U717 ( .A(\rem_74_2/u_div/SumTmp[2][2][3] ), .B(
        \rem_74_2/u_div/SumTmp[6][2][3] ), .S(n399), .Z(n530) );
  EO1 U718 ( .A(\rem_74_2/u_div/SumTmp[4][2][3] ), .B(n190), .C(n557), .D(n530), .Z(n532) );
  ND2 U719 ( .A(n973), .B(n305), .Z(n531) );
  MUX21L U720 ( .A(\rem_74_2/u_div/SumTmp[3][2][2] ), .B(
        \rem_74_2/u_div/SumTmp[7][2][2] ), .S(n399), .Z(n533) );
  EO1 U721 ( .A(\rem_74_2/u_div/SumTmp[5][2][2] ), .B(n302), .C(n557), .D(n533), .Z(n535) );
  ND2 U722 ( .A(\rem_74_2/u_div/SumTmp[1][2][2] ), .B(n305), .Z(n534) );
  ND2 U723 ( .A(n535), .B(n534), .Z(n536) );
  IVA U724 ( .A(n536), .Z(n564) );
  MUX21L U725 ( .A(\rem_74_2/u_div/SumTmp[2][2][2] ), .B(
        \rem_74_2/u_div/SumTmp[6][2][2] ), .S(n79), .Z(n537) );
  EO1 U726 ( .A(\rem_74_2/u_div/SumTmp[4][2][2] ), .B(n302), .C(n557), .D(n537), .Z(n539) );
  ND2 U727 ( .A(n305), .B(input_no[8]), .Z(n538) );
  ND2 U728 ( .A(n539), .B(n538), .Z(n540) );
  IVA U729 ( .A(n540), .Z(n563) );
  MUX21L U730 ( .A(\rem_74_2/u_div/SumTmp[3][2][1] ), .B(
        \rem_74_2/u_div/SumTmp[7][2][1] ), .S(n79), .Z(n541) );
  EO1 U731 ( .A(\rem_74_2/u_div/SumTmp[1][2][1] ), .B(n189), .C(n541), .D(n557), .Z(n543) );
  ND2 U732 ( .A(\rem_74_2/u_div/SumTmp[5][2][1] ), .B(n302), .Z(n542) );
  ND2 U733 ( .A(n543), .B(n542), .Z(n544) );
  MUX21L U734 ( .A(\rem_74_2/u_div/SumTmp[2][2][1] ), .B(
        \rem_74_2/u_div/SumTmp[6][2][1] ), .S(n79), .Z(n545) );
  EO1 U735 ( .A(n189), .B(input_no[7]), .C(n545), .D(n557), .Z(n547) );
  ND2 U736 ( .A(\rem_74_2/u_div/SumTmp[4][2][1] ), .B(n190), .Z(n546) );
  ND2 U737 ( .A(n547), .B(n546), .Z(n548) );
  MUX21L U738 ( .A(\rem_74_2/u_div/SumTmp[3][2][0] ), .B(
        \rem_74_2/u_div/SumTmp[7][2][0] ), .S(n212), .Z(n554) );
  MUX21L U739 ( .A(\rem_74_2/u_div/SumTmp[2][2][0] ), .B(
        \rem_74_2/u_div/SumTmp[6][2][0] ), .S(n212), .Z(n558) );
  MUX21H U740 ( .A(\rem_74_2/u_div/SumTmp[3][1][8] ), .B(
        \rem_74_2/u_div/SumTmp[7][1][8] ), .S(n161), .Z(n570) );
  IVA U741 ( .A(n972), .Z(n572) );
  MUX21L U742 ( .A(\rem_74_2/u_div/SumTmp[2][1][8] ), .B(
        \rem_74_2/u_div/SumTmp[6][1][8] ), .S(n103), .Z(n571) );
  AO4 U743 ( .A(n572), .B(n228), .C(n295), .D(n571), .Z(n573) );
  MUX21H U744 ( .A(\rem_74_2/u_div/SumTmp[3][1][7] ), .B(
        \rem_74_2/u_div/SumTmp[7][1][7] ), .S(n161), .Z(n584) );
  AO11 U745 ( .A(\rem_74_2/u_div/SumTmp[1][1][7] ), .B(n105), .C(n584), .D(
        n246), .E(\rem_74_2/u_div/SumTmp[5][1][7] ), .F(n338), .Z(n589) );
  IVA U746 ( .A(n971), .Z(n586) );
  MUX21L U747 ( .A(\rem_74_2/u_div/SumTmp[2][1][7] ), .B(
        \rem_74_2/u_div/SumTmp[6][1][7] ), .S(n103), .Z(n585) );
  AO4 U748 ( .A(n586), .B(n228), .C(n295), .D(n585), .Z(n587) );
  ND2 U749 ( .A(\rem_74_2/u_div/SumTmp[5][1][6] ), .B(n338), .Z(n590) );
  ND2 U750 ( .A(n628), .B(n968), .Z(n592) );
  MUX21L U751 ( .A(\rem_74_2/u_div/SumTmp[3][1][5] ), .B(
        \rem_74_2/u_div/SumTmp[7][1][5] ), .S(n103), .Z(n594) );
  EO1 U752 ( .A(\rem_74_2/u_div/SumTmp[1][1][5] ), .B(n628), .C(n594), .D(n295), .Z(n596) );
  ND2 U753 ( .A(\rem_74_2/u_div/SumTmp[5][1][5] ), .B(n338), .Z(n595) );
  ND2 U754 ( .A(n596), .B(n595), .Z(n597) );
  MUX21L U755 ( .A(\rem_74_2/u_div/SumTmp[2][1][5] ), .B(
        \rem_74_2/u_div/SumTmp[6][1][5] ), .S(n103), .Z(n598) );
  EO1 U756 ( .A(\rem_74_2/u_div/SumTmp[4][1][5] ), .B(n297), .C(n598), .D(n295), .Z(n600) );
  ND2 U757 ( .A(n628), .B(n967), .Z(n599) );
  ND2 U758 ( .A(n600), .B(n599), .Z(n601) );
  MUX21L U759 ( .A(\rem_74_2/u_div/SumTmp[3][1][4] ), .B(
        \rem_74_2/u_div/SumTmp[7][1][4] ), .S(n104), .Z(n602) );
  EO1 U760 ( .A(\rem_74_2/u_div/SumTmp[1][1][4] ), .B(n227), .C(n602), .D(n630), .Z(n604) );
  ND2 U761 ( .A(\rem_74_2/u_div/SumTmp[5][1][4] ), .B(n338), .Z(n603) );
  MUX21L U762 ( .A(\rem_74_2/u_div/SumTmp[2][1][4] ), .B(
        \rem_74_2/u_div/SumTmp[6][1][4] ), .S(n425), .Z(n605) );
  EO1 U763 ( .A(n227), .B(n964), .C(n605), .D(n630), .Z(n607) );
  ND2 U764 ( .A(\rem_74_2/u_div/SumTmp[4][1][4] ), .B(n338), .Z(n606) );
  MUX21H U765 ( .A(\rem_74_2/u_div/SumTmp[3][1][3] ), .B(
        \rem_74_2/u_div/SumTmp[7][1][3] ), .S(n103), .Z(n608) );
  AO11 U766 ( .A(n246), .B(n608), .C(\rem_74_2/u_div/SumTmp[1][1][3] ), .D(
        n628), .E(\rem_74_2/u_div/SumTmp[5][1][3] ), .F(n338), .Z(n615) );
  MUX21L U767 ( .A(\rem_74_2/u_div/SumTmp[2][1][3] ), .B(
        \rem_74_2/u_div/SumTmp[6][1][3] ), .S(n425), .Z(n610) );
  AO4 U768 ( .A(n610), .B(n630), .C(n609), .D(n629), .Z(n611) );
  MUX21H U769 ( .A(\rem_74_2/u_div/SumTmp[3][1][2] ), .B(
        \rem_74_2/u_div/SumTmp[7][1][2] ), .S(n425), .Z(n616) );
  MUX21L U770 ( .A(\rem_74_2/u_div/SumTmp[2][1][2] ), .B(
        \rem_74_2/u_div/SumTmp[6][1][2] ), .S(n425), .Z(n617) );
  AO4 U771 ( .A(n617), .B(n630), .C(n982), .D(n629), .Z(n618) );
  MUX21H U772 ( .A(\rem_74_2/u_div/SumTmp[3][1][1] ), .B(
        \rem_74_2/u_div/SumTmp[7][1][1] ), .S(n425), .Z(n621) );
  AO11 U773 ( .A(\rem_74_2/u_div/SumTmp[5][1][1] ), .B(n338), .C(
        \rem_74_2/u_div/SumTmp[1][1][1] ), .D(n628), .E(n246), .F(n621), .Z(
        n626) );
  MUX21L U774 ( .A(\rem_74_2/u_div/SumTmp[2][1][1] ), .B(
        \rem_74_2/u_div/SumTmp[6][1][1] ), .S(n424), .Z(n623) );
  AO4 U775 ( .A(n623), .B(n630), .C(n622), .D(n629), .Z(n624) );
  MUX21H U776 ( .A(\rem_74_2/u_div/SumTmp[3][1][0] ), .B(
        \rem_74_2/u_div/SumTmp[7][1][0] ), .S(n425), .Z(n627) );
  AO11 U777 ( .A(\rem_74_2/u_div/SumTmp[5][1][0] ), .B(n297), .C(
        \rem_74_2/u_div/SumTmp[1][1][0] ), .D(n628), .E(n246), .F(n627), .Z(
        n634) );
  MUX21L U778 ( .A(\rem_74_2/u_div/SumTmp[2][1][0] ), .B(
        \rem_74_2/u_div/SumTmp[6][1][0] ), .S(n103), .Z(n631) );
  AO4 U779 ( .A(n631), .B(n630), .C(n433), .D(n629), .Z(n632) );
  MUX21L U780 ( .A(\rem_74/u_div/SumTmp[3][2][5] ), .B(
        \rem_74/u_div/SumTmp[7][2][5] ), .S(n233), .Z(n641) );
  EO1 U781 ( .A(\rem_74/u_div/SumTmp[5][2][5] ), .B(n343), .C(n686), .D(n641), 
        .Z(n643) );
  ND2 U782 ( .A(\rem_74/u_div/SumTmp[1][2][5] ), .B(n364), .Z(n642) );
  MUX21L U783 ( .A(\rem_74/u_div/SumTmp[2][2][5] ), .B(
        \rem_74/u_div/SumTmp[6][2][5] ), .S(n64), .Z(n644) );
  EO1 U784 ( .A(\rem_74/u_div/SumTmp[4][2][5] ), .B(n343), .C(n686), .D(n644), 
        .Z(n646) );
  ND2 U785 ( .A(n949), .B(n364), .Z(n645) );
  MUX21L U786 ( .A(\rem_74/u_div/SumTmp[3][2][4] ), .B(
        \rem_74/u_div/SumTmp[7][2][4] ), .S(n64), .Z(n647) );
  EO1 U787 ( .A(\rem_74/u_div/SumTmp[5][2][4] ), .B(n343), .C(n686), .D(n647), 
        .Z(n649) );
  ND2 U788 ( .A(\rem_74/u_div/SumTmp[1][2][4] ), .B(n364), .Z(n648) );
  MUX21L U789 ( .A(\rem_74/u_div/SumTmp[2][2][4] ), .B(
        \rem_74/u_div/SumTmp[6][2][4] ), .S(n64), .Z(n650) );
  EO1 U790 ( .A(\rem_74/u_div/SumTmp[4][2][4] ), .B(n343), .C(n686), .D(n650), 
        .Z(n652) );
  ND2 U791 ( .A(n948), .B(n364), .Z(n651) );
  MUX21L U792 ( .A(\rem_74/u_div/SumTmp[2][2][3] ), .B(
        \rem_74/u_div/SumTmp[6][2][3] ), .S(n265), .Z(n653) );
  AO4 U793 ( .A(n676), .B(n654), .C(n310), .D(n653), .Z(n656) );
  OR2 U794 ( .A(n656), .B(n118), .Z(n694) );
  MUX21L U795 ( .A(\rem_74/u_div/SumTmp[3][2][3] ), .B(
        \rem_74/u_div/SumTmp[7][2][3] ), .S(n265), .Z(n657) );
  AO4 U796 ( .A(n676), .B(n658), .C(n686), .D(n657), .Z(n659) );
  OR2 U797 ( .A(n116), .B(n659), .Z(n693) );
  AO2 U798 ( .A(\rem_74/u_div/SumTmp[4][2][2] ), .B(n64), .C(input_no[8]), .D(
        n280), .Z(n662) );
  MUX21L U799 ( .A(\rem_74/u_div/SumTmp[2][2][2] ), .B(
        \rem_74/u_div/SumTmp[6][2][2] ), .S(n64), .Z(n661) );
  AO4 U800 ( .A(n676), .B(n662), .C(n686), .D(n661), .Z(n666) );
  AO2 U801 ( .A(\rem_74/u_div/SumTmp[5][2][2] ), .B(n265), .C(
        \rem_74/u_div/SumTmp[1][2][2] ), .D(n280), .Z(n664) );
  MUX21L U802 ( .A(\rem_74/u_div/SumTmp[3][2][2] ), .B(
        \rem_74/u_div/SumTmp[7][2][2] ), .S(n265), .Z(n663) );
  AO4 U803 ( .A(n676), .B(n664), .C(n686), .D(n663), .Z(n665) );
  AO2 U804 ( .A(\rem_74/u_div/SumTmp[4][2][1] ), .B(n64), .C(input_no[7]), .D(
        n280), .Z(n669) );
  MUX21L U805 ( .A(\rem_74/u_div/SumTmp[2][2][1] ), .B(
        \rem_74/u_div/SumTmp[6][2][1] ), .S(n265), .Z(n668) );
  AO4 U806 ( .A(n309), .B(n669), .C(n668), .D(n310), .Z(n673) );
  MUX21L U807 ( .A(\rem_74/u_div/SumTmp[3][2][1] ), .B(
        \rem_74/u_div/SumTmp[7][2][1] ), .S(n64), .Z(n677) );
  AO2 U808 ( .A(\rem_74/u_div/SumTmp[5][2][1] ), .B(n64), .C(
        \rem_74/u_div/SumTmp[1][2][1] ), .D(n280), .Z(n675) );
  AO4 U809 ( .A(n677), .B(n686), .C(n309), .D(n675), .Z(n678) );
  AO2 U810 ( .A(\rem_74/u_div/SumTmp[5][2][0] ), .B(n265), .C(
        \rem_74/u_div/SumTmp[1][2][0] ), .D(n280), .Z(n680) );
  AO2 U811 ( .A(\rem_74/u_div/SumTmp[4][2][0] ), .B(n64), .C(input_no[6]), .D(
        n280), .Z(n681) );
  MUX21L U812 ( .A(\rem_74/u_div/SumTmp[3][2][0] ), .B(
        \rem_74/u_div/SumTmp[7][2][0] ), .S(n265), .Z(n685) );
  MUX21L U813 ( .A(\rem_74/u_div/SumTmp[2][2][0] ), .B(
        \rem_74/u_div/SumTmp[6][2][0] ), .S(n64), .Z(n683) );
  AN2P U814 ( .A(n694), .B(n693), .Z(n943) );
  ND2 U815 ( .A(n235), .B(n293), .Z(n709) );
  IVA U816 ( .A(n709), .Z(n739) );
  MUX21H U817 ( .A(\rem_74/u_div/SumTmp[3][1][8] ), .B(
        \rem_74/u_div/SumTmp[7][1][8] ), .S(n164), .Z(n695) );
  AO11 U818 ( .A(\rem_74/u_div/SumTmp[1][1][8] ), .B(n739), .C(n695), .D(n230), 
        .E(\rem_74/u_div/SumTmp[5][1][8] ), .F(n173), .Z(n706) );
  IVA U819 ( .A(n946), .Z(n697) );
  MUX21L U820 ( .A(\rem_74/u_div/SumTmp[2][1][8] ), .B(
        \rem_74/u_div/SumTmp[6][1][8] ), .S(n66), .Z(n696) );
  AO4 U821 ( .A(n697), .B(n709), .C(n769), .D(n696), .Z(n698) );
  AN3 U822 ( .A(\rem_74/u_div/CryOut[1][1] ), .B(n235), .C(n293), .Z(n703) );
  MUX21H U823 ( .A(\rem_74/u_div/SumTmp[3][1][7] ), .B(
        \rem_74/u_div/SumTmp[7][1][7] ), .S(n311), .Z(n707) );
  AO11 U824 ( .A(\rem_74/u_div/SumTmp[1][1][7] ), .B(n739), .C(n707), .D(n230), 
        .E(\rem_74/u_div/SumTmp[5][1][7] ), .F(n173), .Z(n713) );
  IVA U825 ( .A(n332), .Z(n710) );
  MUX21L U826 ( .A(\rem_74/u_div/SumTmp[2][1][7] ), .B(
        \rem_74/u_div/SumTmp[6][1][7] ), .S(n66), .Z(n708) );
  AO4 U827 ( .A(n710), .B(n709), .C(n769), .D(n708), .Z(n711) );
  MUX21L U828 ( .A(\rem_74/u_div/SumTmp[3][1][6] ), .B(
        \rem_74/u_div/SumTmp[7][1][6] ), .S(n422), .Z(n714) );
  AN3 U829 ( .A(\rem_74/u_div/SumTmp[1][1][6] ), .B(n357), .C(n769), .Z(n715)
         );
  AO1P U830 ( .A(\rem_74/u_div/SumTmp[5][1][6] ), .B(n339), .C(n716), .D(n715), 
        .Z(n721) );
  AN3 U831 ( .A(n216), .B(n357), .C(n769), .Z(n719) );
  MUX21L U832 ( .A(\rem_74/u_div/SumTmp[2][1][6] ), .B(
        \rem_74/u_div/SumTmp[6][1][6] ), .S(n422), .Z(n717) );
  AO1P U833 ( .A(\rem_74/u_div/SumTmp[4][1][6] ), .B(n339), .C(n719), .D(n718), 
        .Z(n720) );
  MUX21L U834 ( .A(\rem_74/u_div/SumTmp[3][1][5] ), .B(
        \rem_74/u_div/SumTmp[7][1][5] ), .S(n422), .Z(n722) );
  AN3 U835 ( .A(\rem_74/u_div/SumTmp[1][1][5] ), .B(n356), .C(n753), .Z(n723)
         );
  AO1P U836 ( .A(\rem_74/u_div/SumTmp[5][1][5] ), .B(n173), .C(n724), .D(n723), 
        .Z(n729) );
  AN3 U837 ( .A(n291), .B(n158), .C(n753), .Z(n727) );
  MUX21L U838 ( .A(\rem_74/u_div/SumTmp[2][1][5] ), .B(
        \rem_74/u_div/SumTmp[6][1][5] ), .S(n358), .Z(n725) );
  AO1P U839 ( .A(\rem_74/u_div/SumTmp[4][1][5] ), .B(n173), .C(n727), .D(n726), 
        .Z(n728) );
  AO2 U840 ( .A(\rem_74/u_div/SumTmp[4][1][4] ), .B(n422), .C(n211), .D(n158), 
        .Z(n731) );
  MUX21L U841 ( .A(\rem_74/u_div/SumTmp[2][1][4] ), .B(
        \rem_74/u_div/SumTmp[6][1][4] ), .S(n359), .Z(n730) );
  AO4 U842 ( .A(n172), .B(n731), .C(n730), .D(n180), .Z(n735) );
  AO2 U843 ( .A(\rem_74/u_div/SumTmp[5][1][4] ), .B(n66), .C(
        \rem_74/u_div/SumTmp[1][1][4] ), .D(n357), .Z(n733) );
  MUX21L U844 ( .A(\rem_74/u_div/SumTmp[3][1][4] ), .B(
        \rem_74/u_div/SumTmp[7][1][4] ), .S(n164), .Z(n732) );
  AO4 U845 ( .A(n172), .B(n733), .C(n732), .D(n180), .Z(n734) );
  MUX21L U846 ( .A(\rem_74/u_div/SumTmp[3][1][3] ), .B(
        \rem_74/u_div/SumTmp[7][1][3] ), .S(n164), .Z(n738) );
  AO2 U847 ( .A(\rem_74/u_div/SumTmp[1][1][3] ), .B(n739), .C(
        \rem_74/u_div/SumTmp[5][1][3] ), .D(n339), .Z(n737) );
  MUX21L U848 ( .A(\rem_74/u_div/SumTmp[2][1][3] ), .B(
        \rem_74/u_div/SumTmp[6][1][3] ), .S(n311), .Z(n741) );
  AO2 U849 ( .A(n174), .B(n739), .C(\rem_74/u_div/SumTmp[4][1][3] ), .D(n339), 
        .Z(n740) );
  AO2 U850 ( .A(\rem_74/u_div/SumTmp[4][1][2] ), .B(n422), .C(input_no[5]), 
        .D(n357), .Z(n745) );
  MUX21L U851 ( .A(\rem_74/u_div/SumTmp[2][1][2] ), .B(
        \rem_74/u_div/SumTmp[6][1][2] ), .S(n359), .Z(n744) );
  AO4 U852 ( .A(n172), .B(n745), .C(n744), .D(n753), .Z(n749) );
  AO2 U853 ( .A(\rem_74/u_div/SumTmp[5][1][2] ), .B(n422), .C(
        \rem_74/u_div/SumTmp[1][1][2] ), .D(n357), .Z(n747) );
  MUX21L U854 ( .A(\rem_74/u_div/SumTmp[3][1][2] ), .B(
        \rem_74/u_div/SumTmp[7][1][2] ), .S(n359), .Z(n746) );
  AO4 U855 ( .A(n172), .B(n747), .C(n746), .D(n753), .Z(n748) );
  AO2 U856 ( .A(\rem_74/u_div/SumTmp[4][1][1] ), .B(n422), .C(input_no[4]), 
        .D(n357), .Z(n752) );
  MUX21L U857 ( .A(\rem_74/u_div/SumTmp[2][1][1] ), .B(
        \rem_74/u_div/SumTmp[6][1][1] ), .S(n66), .Z(n751) );
  AO4 U858 ( .A(n172), .B(n752), .C(n751), .D(n180), .Z(n758) );
  AO2 U859 ( .A(\rem_74/u_div/SumTmp[5][1][1] ), .B(n422), .C(
        \rem_74/u_div/SumTmp[1][1][1] ), .D(n356), .Z(n755) );
  MUX21L U860 ( .A(\rem_74/u_div/SumTmp[3][1][1] ), .B(
        \rem_74/u_div/SumTmp[7][1][1] ), .S(n66), .Z(n754) );
  AO4 U861 ( .A(n172), .B(n755), .C(n754), .D(n180), .Z(n756) );
  MUX21L U862 ( .A(\rem_74/u_div/SumTmp[3][1][0] ), .B(
        \rem_74/u_div/SumTmp[7][1][0] ), .S(n359), .Z(n763) );
  MUX21L U863 ( .A(\rem_74/u_div/CryOut[3][1] ), .B(n234), .S(n358), .Z(n760)
         );
  IVA U864 ( .A(n760), .Z(n762) );
  MUX21L U865 ( .A(\rem_74/u_div/SumTmp[2][1][0] ), .B(
        \rem_74/u_div/SumTmp[6][1][0] ), .S(n359), .Z(n761) );
  AO2 U866 ( .A(\rem_74/u_div/SumTmp[4][1][0] ), .B(n422), .C(input_no[3]), 
        .D(n357), .Z(n767) );
  AO4 U867 ( .A(\rem_74/u_div/CryOut[1][1] ), .B(n423), .C(
        \rem_74/u_div/CryOut[5][1] ), .D(n293), .Z(n766) );
  AO2 U868 ( .A(\rem_74/u_div/SumTmp[5][1][0] ), .B(n422), .C(
        \rem_74/u_div/SumTmp[1][1][0] ), .D(n357), .Z(n765) );
  AO2 U869 ( .A(n767), .B(n766), .C(n765), .D(n764), .Z(n768) );
  MUX21L U870 ( .A(\rem_74/u_div/SumTmp[3][0][5] ), .B(
        \rem_74/u_div/SumTmp[7][0][5] ), .S(n315), .Z(n772) );
  EO1 U871 ( .A(\rem_74/u_div/SumTmp[1][0][5] ), .B(n342), .C(n772), .D(n253), 
        .Z(n775) );
  ND2 U872 ( .A(\rem_74/u_div/SumTmp[5][0][5] ), .B(n155), .Z(n774) );
  ND2 U873 ( .A(n775), .B(n774), .Z(n784) );
  MUX21L U874 ( .A(\rem_74/u_div/SumTmp[2][0][5] ), .B(
        \rem_74/u_div/SumTmp[6][0][5] ), .S(n68), .Z(n776) );
  EON1 U875 ( .A(n776), .B(n828), .C(\rem_74/u_div/SumTmp[4][0][5] ), .D(n152), 
        .Z(n783) );
  MUX21L U876 ( .A(\rem_74/u_div/CryOut[3][0] ), .B(
        \rem_74/u_div/CryOut[7][0] ), .S(n162), .Z(n781) );
  AO2 U877 ( .A(\rem_74/u_div/CryOut[6][0] ), .B(\rem_74/quotient[2] ), .C(
        \rem_74/u_div/CryOut[2][0] ), .D(n312), .Z(n780) );
  ND3 U878 ( .A(\rem_74/u_div/CryOut[1][0] ), .B(n163), .C(n777), .Z(n779) );
  MUX21L U879 ( .A(\rem_74/u_div/SumTmp[3][0][4] ), .B(
        \rem_74/u_div/SumTmp[7][0][4] ), .S(n315), .Z(n785) );
  EO1 U880 ( .A(\rem_74/u_div/SumTmp[1][0][4] ), .B(n342), .C(n785), .D(n253), 
        .Z(n787) );
  ND2 U881 ( .A(\rem_74/u_div/SumTmp[5][0][4] ), .B(n156), .Z(n786) );
  ND2 U882 ( .A(n787), .B(n786), .Z(n790) );
  MUX21L U883 ( .A(\rem_74/u_div/SumTmp[2][0][4] ), .B(
        \rem_74/u_div/SumTmp[6][0][4] ), .S(n315), .Z(n788) );
  EON1 U884 ( .A(n788), .B(n828), .C(\rem_74/u_div/SumTmp[4][0][4] ), .D(n152), 
        .Z(n789) );
  MUX21H U885 ( .A(\rem_74/u_div/SumTmp[3][0][1] ), .B(
        \rem_74/u_div/SumTmp[7][0][1] ), .S(n298), .Z(n793) );
  AO11 U886 ( .A(\rem_74/u_div/SumTmp[5][0][1] ), .B(n156), .C(n793), .D(n827), 
        .E(\rem_74/u_div/SumTmp[1][0][1] ), .F(n342), .Z(n796) );
  MUX21L U887 ( .A(\rem_74/u_div/SumTmp[2][0][1] ), .B(
        \rem_74/u_div/SumTmp[6][0][1] ), .S(n315), .Z(n794) );
  EO1 U888 ( .A(\rem_74/u_div/SumTmp[4][0][1] ), .B(n152), .C(n828), .D(n794), 
        .Z(n795) );
  MUX21H U889 ( .A(\rem_74/u_div/SumTmp[3][0][9] ), .B(
        \rem_74/u_div/SumTmp[7][0][9] ), .S(n315), .Z(n797) );
  AO11 U890 ( .A(n827), .B(n797), .C(\rem_74/u_div/SumTmp[1][0][9] ), .D(n342), 
        .E(\rem_74/u_div/SumTmp[5][0][9] ), .F(n154), .Z(n801) );
  AN3 U891 ( .A(\rem_74/u_div/SumTmp[6][0][9] ), .B(n298), .C(n70), .Z(n799)
         );
  MUX21H U892 ( .A(\rem_74/u_div/SumTmp[3][0][0] ), .B(
        \rem_74/u_div/SumTmp[7][0][0] ), .S(n298), .Z(n802) );
  AO11 U893 ( .A(\rem_74/u_div/SumTmp[5][0][0] ), .B(n155), .C(n802), .D(n827), 
        .E(\rem_74/u_div/SumTmp[1][0][0] ), .F(n342), .Z(n806) );
  NR2P U894 ( .A(n828), .B(n803), .Z(n804) );
  AO1P U895 ( .A(\rem_74/u_div/SumTmp[4][0][0] ), .B(n155), .C(n342), .D(n804), 
        .Z(n805) );
  AO11 U896 ( .A(n827), .B(n807), .C(\rem_74/u_div/SumTmp[1][0][3] ), .D(n342), 
        .E(\rem_74/u_div/SumTmp[5][0][3] ), .F(n151), .Z(n810) );
  MUX21L U897 ( .A(\rem_74/u_div/SumTmp[2][0][3] ), .B(
        \rem_74/u_div/SumTmp[6][0][3] ), .S(n315), .Z(n808) );
  EO1 U898 ( .A(\rem_74/u_div/SumTmp[4][0][3] ), .B(n152), .C(n808), .D(n828), 
        .Z(n809) );
  AO11 U899 ( .A(\rem_74/u_div/SumTmp[5][0][2] ), .B(n151), .C(n814), .D(n827), 
        .E(\rem_74/u_div/SumTmp[1][0][2] ), .F(n342), .Z(n817) );
  MUX21L U900 ( .A(\rem_74/u_div/SumTmp[2][0][2] ), .B(
        \rem_74/u_div/SumTmp[6][0][2] ), .S(n315), .Z(n815) );
  EO1 U901 ( .A(\rem_74/u_div/SumTmp[4][0][2] ), .B(n154), .C(n828), .D(n815), 
        .Z(n816) );
  AO11 U902 ( .A(n827), .B(n818), .C(\rem_74/u_div/SumTmp[1][0][8] ), .D(n342), 
        .E(\rem_74/u_div/SumTmp[5][0][8] ), .F(n156), .Z(n821) );
  MUX21L U903 ( .A(\rem_74/u_div/SumTmp[2][0][8] ), .B(
        \rem_74/u_div/SumTmp[6][0][8] ), .S(n315), .Z(n819) );
  EO1 U904 ( .A(\rem_74/u_div/SumTmp[4][0][8] ), .B(n153), .C(n819), .D(n828), 
        .Z(n820) );
  MUX21H U905 ( .A(\rem_74/u_div/SumTmp[3][0][7] ), .B(
        \rem_74/u_div/SumTmp[7][0][7] ), .S(n315), .Z(n822) );
  AO11 U906 ( .A(n827), .B(n822), .C(\rem_74/u_div/SumTmp[1][0][7] ), .D(n342), 
        .E(\rem_74/u_div/SumTmp[5][0][7] ), .F(n153), .Z(n825) );
  MUX21L U907 ( .A(\rem_74/u_div/SumTmp[2][0][7] ), .B(
        \rem_74/u_div/SumTmp[6][0][7] ), .S(n315), .Z(n823) );
  EO1 U908 ( .A(\rem_74/u_div/SumTmp[4][0][7] ), .B(n154), .C(n823), .D(n828), 
        .Z(n824) );
  MUX21H U909 ( .A(\rem_74/u_div/SumTmp[3][0][6] ), .B(
        \rem_74/u_div/SumTmp[7][0][6] ), .S(n315), .Z(n826) );
  AO11 U910 ( .A(n827), .B(n826), .C(\rem_74/u_div/SumTmp[1][0][6] ), .D(n342), 
        .E(\rem_74/u_div/SumTmp[5][0][6] ), .F(n154), .Z(n832) );
  MUX21L U911 ( .A(\rem_74/u_div/SumTmp[2][0][6] ), .B(
        \rem_74/u_div/SumTmp[6][0][6] ), .S(n315), .Z(n829) );
  EO1 U912 ( .A(\rem_74/u_div/SumTmp[4][0][6] ), .B(n154), .C(n829), .D(n828), 
        .Z(n831) );
  OR3 U913 ( .A(n923), .B(n836), .C(n835), .Z(n892) );
  MUX21L U914 ( .A(n106), .B(n109), .S(n72), .Z(n907) );
  NR5 U915 ( .A(\rem_74_2/u_div/SumTmp[2][0][9] ), .B(
        \rem_74_2/u_div/SumTmp[2][0][2] ), .C(\rem_74_2/u_div/SumTmp[2][0][3] ), .D(\rem_74_2/u_div/SumTmp[2][0][4] ), .E(\rem_74_2/u_div/SumTmp[2][0][5] ), 
        .Z(n909) );
  OR3 U916 ( .A(\rem_74_2/u_div/SumTmp[4][0][1] ), .B(
        \rem_74_2/u_div/SumTmp[4][0][2] ), .C(\rem_74_2/u_div/SumTmp[4][0][5] ), .Z(n893) );
  OR3 U917 ( .A(\rem_74_2/u_div/SumTmp[4][0][7] ), .B(n109), .C(n893), .Z(n894) );
  ND2 U918 ( .A(n895), .B(n894), .Z(n908) );
  OR3 U919 ( .A(\rem_74_2/u_div/SumTmp[2][0][0] ), .B(\rem_74_2/quotient[2] ), 
        .C(\rem_74_2/u_div/SumTmp[2][0][7] ), .Z(n897) );
  OR3 U920 ( .A(\rem_74_2/u_div/SumTmp[6][0][0] ), .B(n119), .C(
        \rem_74_2/u_div/SumTmp[6][0][7] ), .Z(n896) );
  ND2 U921 ( .A(n897), .B(n896), .Z(n906) );
  OR3 U922 ( .A(\rem_74_2/u_div/SumTmp[6][0][1] ), .B(
        \rem_74_2/u_div/SumTmp[6][0][6] ), .C(\rem_74_2/u_div/CryOut[7][0] ), 
        .Z(n903) );
  OR3 U923 ( .A(\rem_74_2/u_div/SumTmp[2][0][1] ), .B(
        \rem_74_2/u_div/SumTmp[2][0][6] ), .C(\rem_74_2/u_div/CryOut[3][0] ), 
        .Z(n901) );
  ND2 U924 ( .A(input_no[1]), .B(\state[0] ), .Z(n911) );
  AO4 U925 ( .A(n913), .B(n912), .C(n911), .D(n910), .Z(n919) );
  IVA U926 ( .A(n919), .Z(n927) );
  ND2 U927 ( .A(n915), .B(n914), .Z(n926) );
  ND3 U928 ( .A(n336), .B(n341), .C(n346), .Z(n922) );
  NR8P U929 ( .A(n923), .B(n922), .C(n921), .D(n920), .E(n919), .F(n918), .G(
        n917), .H(n916), .Z(n924) );
  AO1P U930 ( .A(n927), .B(n926), .C(n925), .D(n924), .Z(n58) );
  NR2 U935 ( .A(input_no[1]), .B(input_no[0]), .Z(n981) );
endmodule

